-----------------------------------------------------------------------------
--! @file
--! @copyright Copyright 2015 GNSS Sensor Ltd. All right reserved.
--! @author    Sergey Khabarov - sergeykhbr@gmail.com
--! @brief     Matrix correlator 4096 samples length
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
library commonlib;
use commonlib.types_common.all;
library gnsslib;
use gnsslib.types_fse_v2.all;

entity Matrix24 is
port (
    i_nrst          : in std_logic;
    i_clk           : in std_logic;
    i_ena           : in std_logic;
    i_re_im         : in std_logic;
    i_prn           : in std_logic_vector(1024-1 downto 0);
    i_I             : in std_logic_vector(2*1024-1 downto 0);
    i_Q             : in std_logic_vector(2*1024-1 downto 0);
    o_lvl1          : out std_logic_vector(512*4-1 downto 0)
);
end;

architecture rtl of Matrix24 is


type regtype is record
  Lvl1     : std_logic_vector(512*4-1 downto 0);
end record;

signal r, rin : regtype;

begin

  comb : process (r, i_nrst, i_ena, i_re_im, i_prn, i_I, i_Q)
  variable v : regtype;
  variable wbPartMux : std_logic_vector(2*1024-1 downto 0);
  variable wbMult : std_logic_vector(3*1024-1 downto 0);
  
  begin
    
    --v := r;

    if i_re_im = '1' then 
      wbPartMux := i_Q;
    else
      wbPartMux := i_I;
    end if;
    
    wbMult(2 downto 0) := (wbPartMux(1) xor i_prn(0)) & (not wbPartMux(0) xor i_prn(0)) & '1';
    wbMult(5 downto 3) := (wbPartMux(3) xor i_prn(1)) & (not wbPartMux(2) xor i_prn(1)) & '1';
    wbMult(8 downto 6) := (wbPartMux(5) xor i_prn(2)) & (not wbPartMux(4) xor i_prn(2)) & '1';
    wbMult(11 downto 9) := (wbPartMux(7) xor i_prn(3)) & (not wbPartMux(6) xor i_prn(3)) & '1';
    wbMult(14 downto 12) := (wbPartMux(9) xor i_prn(4)) & (not wbPartMux(8) xor i_prn(4)) & '1';
    wbMult(17 downto 15) := (wbPartMux(11) xor i_prn(5)) & (not wbPartMux(10) xor i_prn(5)) & '1';
    wbMult(20 downto 18) := (wbPartMux(13) xor i_prn(6)) & (not wbPartMux(12) xor i_prn(6)) & '1';
    wbMult(23 downto 21) := (wbPartMux(15) xor i_prn(7)) & (not wbPartMux(14) xor i_prn(7)) & '1';
    wbMult(26 downto 24) := (wbPartMux(17) xor i_prn(8)) & (not wbPartMux(16) xor i_prn(8)) & '1';
    wbMult(29 downto 27) := (wbPartMux(19) xor i_prn(9)) & (not wbPartMux(18) xor i_prn(9)) & '1';
    wbMult(32 downto 30) := (wbPartMux(21) xor i_prn(10)) & (not wbPartMux(20) xor i_prn(10)) & '1';
    wbMult(35 downto 33) := (wbPartMux(23) xor i_prn(11)) & (not wbPartMux(22) xor i_prn(11)) & '1';
    wbMult(38 downto 36) := (wbPartMux(25) xor i_prn(12)) & (not wbPartMux(24) xor i_prn(12)) & '1';
    wbMult(41 downto 39) := (wbPartMux(27) xor i_prn(13)) & (not wbPartMux(26) xor i_prn(13)) & '1';
    wbMult(44 downto 42) := (wbPartMux(29) xor i_prn(14)) & (not wbPartMux(28) xor i_prn(14)) & '1';
    wbMult(47 downto 45) := (wbPartMux(31) xor i_prn(15)) & (not wbPartMux(30) xor i_prn(15)) & '1';
    wbMult(50 downto 48) := (wbPartMux(33) xor i_prn(16)) & (not wbPartMux(32) xor i_prn(16)) & '1';
    wbMult(53 downto 51) := (wbPartMux(35) xor i_prn(17)) & (not wbPartMux(34) xor i_prn(17)) & '1';
    wbMult(56 downto 54) := (wbPartMux(37) xor i_prn(18)) & (not wbPartMux(36) xor i_prn(18)) & '1';
    wbMult(59 downto 57) := (wbPartMux(39) xor i_prn(19)) & (not wbPartMux(38) xor i_prn(19)) & '1';
    wbMult(62 downto 60) := (wbPartMux(41) xor i_prn(20)) & (not wbPartMux(40) xor i_prn(20)) & '1';
    wbMult(65 downto 63) := (wbPartMux(43) xor i_prn(21)) & (not wbPartMux(42) xor i_prn(21)) & '1';
    wbMult(68 downto 66) := (wbPartMux(45) xor i_prn(22)) & (not wbPartMux(44) xor i_prn(22)) & '1';
    wbMult(71 downto 69) := (wbPartMux(47) xor i_prn(23)) & (not wbPartMux(46) xor i_prn(23)) & '1';
    wbMult(74 downto 72) := (wbPartMux(49) xor i_prn(24)) & (not wbPartMux(48) xor i_prn(24)) & '1';
    wbMult(77 downto 75) := (wbPartMux(51) xor i_prn(25)) & (not wbPartMux(50) xor i_prn(25)) & '1';
    wbMult(80 downto 78) := (wbPartMux(53) xor i_prn(26)) & (not wbPartMux(52) xor i_prn(26)) & '1';
    wbMult(83 downto 81) := (wbPartMux(55) xor i_prn(27)) & (not wbPartMux(54) xor i_prn(27)) & '1';
    wbMult(86 downto 84) := (wbPartMux(57) xor i_prn(28)) & (not wbPartMux(56) xor i_prn(28)) & '1';
    wbMult(89 downto 87) := (wbPartMux(59) xor i_prn(29)) & (not wbPartMux(58) xor i_prn(29)) & '1';
    wbMult(92 downto 90) := (wbPartMux(61) xor i_prn(30)) & (not wbPartMux(60) xor i_prn(30)) & '1';
    wbMult(95 downto 93) := (wbPartMux(63) xor i_prn(31)) & (not wbPartMux(62) xor i_prn(31)) & '1';
    wbMult(98 downto 96) := (wbPartMux(65) xor i_prn(32)) & (not wbPartMux(64) xor i_prn(32)) & '1';
    wbMult(101 downto 99) := (wbPartMux(67) xor i_prn(33)) & (not wbPartMux(66) xor i_prn(33)) & '1';
    wbMult(104 downto 102) := (wbPartMux(69) xor i_prn(34)) & (not wbPartMux(68) xor i_prn(34)) & '1';
    wbMult(107 downto 105) := (wbPartMux(71) xor i_prn(35)) & (not wbPartMux(70) xor i_prn(35)) & '1';
    wbMult(110 downto 108) := (wbPartMux(73) xor i_prn(36)) & (not wbPartMux(72) xor i_prn(36)) & '1';
    wbMult(113 downto 111) := (wbPartMux(75) xor i_prn(37)) & (not wbPartMux(74) xor i_prn(37)) & '1';
    wbMult(116 downto 114) := (wbPartMux(77) xor i_prn(38)) & (not wbPartMux(76) xor i_prn(38)) & '1';
    wbMult(119 downto 117) := (wbPartMux(79) xor i_prn(39)) & (not wbPartMux(78) xor i_prn(39)) & '1';
    wbMult(122 downto 120) := (wbPartMux(81) xor i_prn(40)) & (not wbPartMux(80) xor i_prn(40)) & '1';
    wbMult(125 downto 123) := (wbPartMux(83) xor i_prn(41)) & (not wbPartMux(82) xor i_prn(41)) & '1';
    wbMult(128 downto 126) := (wbPartMux(85) xor i_prn(42)) & (not wbPartMux(84) xor i_prn(42)) & '1';
    wbMult(131 downto 129) := (wbPartMux(87) xor i_prn(43)) & (not wbPartMux(86) xor i_prn(43)) & '1';
    wbMult(134 downto 132) := (wbPartMux(89) xor i_prn(44)) & (not wbPartMux(88) xor i_prn(44)) & '1';
    wbMult(137 downto 135) := (wbPartMux(91) xor i_prn(45)) & (not wbPartMux(90) xor i_prn(45)) & '1';
    wbMult(140 downto 138) := (wbPartMux(93) xor i_prn(46)) & (not wbPartMux(92) xor i_prn(46)) & '1';
    wbMult(143 downto 141) := (wbPartMux(95) xor i_prn(47)) & (not wbPartMux(94) xor i_prn(47)) & '1';
    wbMult(146 downto 144) := (wbPartMux(97) xor i_prn(48)) & (not wbPartMux(96) xor i_prn(48)) & '1';
    wbMult(149 downto 147) := (wbPartMux(99) xor i_prn(49)) & (not wbPartMux(98) xor i_prn(49)) & '1';
    wbMult(152 downto 150) := (wbPartMux(101) xor i_prn(50)) & (not wbPartMux(100) xor i_prn(50)) & '1';
    wbMult(155 downto 153) := (wbPartMux(103) xor i_prn(51)) & (not wbPartMux(102) xor i_prn(51)) & '1';
    wbMult(158 downto 156) := (wbPartMux(105) xor i_prn(52)) & (not wbPartMux(104) xor i_prn(52)) & '1';
    wbMult(161 downto 159) := (wbPartMux(107) xor i_prn(53)) & (not wbPartMux(106) xor i_prn(53)) & '1';
    wbMult(164 downto 162) := (wbPartMux(109) xor i_prn(54)) & (not wbPartMux(108) xor i_prn(54)) & '1';
    wbMult(167 downto 165) := (wbPartMux(111) xor i_prn(55)) & (not wbPartMux(110) xor i_prn(55)) & '1';
    wbMult(170 downto 168) := (wbPartMux(113) xor i_prn(56)) & (not wbPartMux(112) xor i_prn(56)) & '1';
    wbMult(173 downto 171) := (wbPartMux(115) xor i_prn(57)) & (not wbPartMux(114) xor i_prn(57)) & '1';
    wbMult(176 downto 174) := (wbPartMux(117) xor i_prn(58)) & (not wbPartMux(116) xor i_prn(58)) & '1';
    wbMult(179 downto 177) := (wbPartMux(119) xor i_prn(59)) & (not wbPartMux(118) xor i_prn(59)) & '1';
    wbMult(182 downto 180) := (wbPartMux(121) xor i_prn(60)) & (not wbPartMux(120) xor i_prn(60)) & '1';
    wbMult(185 downto 183) := (wbPartMux(123) xor i_prn(61)) & (not wbPartMux(122) xor i_prn(61)) & '1';
    wbMult(188 downto 186) := (wbPartMux(125) xor i_prn(62)) & (not wbPartMux(124) xor i_prn(62)) & '1';
    wbMult(191 downto 189) := (wbPartMux(127) xor i_prn(63)) & (not wbPartMux(126) xor i_prn(63)) & '1';
    wbMult(194 downto 192) := (wbPartMux(129) xor i_prn(64)) & (not wbPartMux(128) xor i_prn(64)) & '1';
    wbMult(197 downto 195) := (wbPartMux(131) xor i_prn(65)) & (not wbPartMux(130) xor i_prn(65)) & '1';
    wbMult(200 downto 198) := (wbPartMux(133) xor i_prn(66)) & (not wbPartMux(132) xor i_prn(66)) & '1';
    wbMult(203 downto 201) := (wbPartMux(135) xor i_prn(67)) & (not wbPartMux(134) xor i_prn(67)) & '1';
    wbMult(206 downto 204) := (wbPartMux(137) xor i_prn(68)) & (not wbPartMux(136) xor i_prn(68)) & '1';
    wbMult(209 downto 207) := (wbPartMux(139) xor i_prn(69)) & (not wbPartMux(138) xor i_prn(69)) & '1';
    wbMult(212 downto 210) := (wbPartMux(141) xor i_prn(70)) & (not wbPartMux(140) xor i_prn(70)) & '1';
    wbMult(215 downto 213) := (wbPartMux(143) xor i_prn(71)) & (not wbPartMux(142) xor i_prn(71)) & '1';
    wbMult(218 downto 216) := (wbPartMux(145) xor i_prn(72)) & (not wbPartMux(144) xor i_prn(72)) & '1';
    wbMult(221 downto 219) := (wbPartMux(147) xor i_prn(73)) & (not wbPartMux(146) xor i_prn(73)) & '1';
    wbMult(224 downto 222) := (wbPartMux(149) xor i_prn(74)) & (not wbPartMux(148) xor i_prn(74)) & '1';
    wbMult(227 downto 225) := (wbPartMux(151) xor i_prn(75)) & (not wbPartMux(150) xor i_prn(75)) & '1';
    wbMult(230 downto 228) := (wbPartMux(153) xor i_prn(76)) & (not wbPartMux(152) xor i_prn(76)) & '1';
    wbMult(233 downto 231) := (wbPartMux(155) xor i_prn(77)) & (not wbPartMux(154) xor i_prn(77)) & '1';
    wbMult(236 downto 234) := (wbPartMux(157) xor i_prn(78)) & (not wbPartMux(156) xor i_prn(78)) & '1';
    wbMult(239 downto 237) := (wbPartMux(159) xor i_prn(79)) & (not wbPartMux(158) xor i_prn(79)) & '1';
    wbMult(242 downto 240) := (wbPartMux(161) xor i_prn(80)) & (not wbPartMux(160) xor i_prn(80)) & '1';
    wbMult(245 downto 243) := (wbPartMux(163) xor i_prn(81)) & (not wbPartMux(162) xor i_prn(81)) & '1';
    wbMult(248 downto 246) := (wbPartMux(165) xor i_prn(82)) & (not wbPartMux(164) xor i_prn(82)) & '1';
    wbMult(251 downto 249) := (wbPartMux(167) xor i_prn(83)) & (not wbPartMux(166) xor i_prn(83)) & '1';
    wbMult(254 downto 252) := (wbPartMux(169) xor i_prn(84)) & (not wbPartMux(168) xor i_prn(84)) & '1';
    wbMult(257 downto 255) := (wbPartMux(171) xor i_prn(85)) & (not wbPartMux(170) xor i_prn(85)) & '1';
    wbMult(260 downto 258) := (wbPartMux(173) xor i_prn(86)) & (not wbPartMux(172) xor i_prn(86)) & '1';
    wbMult(263 downto 261) := (wbPartMux(175) xor i_prn(87)) & (not wbPartMux(174) xor i_prn(87)) & '1';
    wbMult(266 downto 264) := (wbPartMux(177) xor i_prn(88)) & (not wbPartMux(176) xor i_prn(88)) & '1';
    wbMult(269 downto 267) := (wbPartMux(179) xor i_prn(89)) & (not wbPartMux(178) xor i_prn(89)) & '1';
    wbMult(272 downto 270) := (wbPartMux(181) xor i_prn(90)) & (not wbPartMux(180) xor i_prn(90)) & '1';
    wbMult(275 downto 273) := (wbPartMux(183) xor i_prn(91)) & (not wbPartMux(182) xor i_prn(91)) & '1';
    wbMult(278 downto 276) := (wbPartMux(185) xor i_prn(92)) & (not wbPartMux(184) xor i_prn(92)) & '1';
    wbMult(281 downto 279) := (wbPartMux(187) xor i_prn(93)) & (not wbPartMux(186) xor i_prn(93)) & '1';
    wbMult(284 downto 282) := (wbPartMux(189) xor i_prn(94)) & (not wbPartMux(188) xor i_prn(94)) & '1';
    wbMult(287 downto 285) := (wbPartMux(191) xor i_prn(95)) & (not wbPartMux(190) xor i_prn(95)) & '1';
    wbMult(290 downto 288) := (wbPartMux(193) xor i_prn(96)) & (not wbPartMux(192) xor i_prn(96)) & '1';
    wbMult(293 downto 291) := (wbPartMux(195) xor i_prn(97)) & (not wbPartMux(194) xor i_prn(97)) & '1';
    wbMult(296 downto 294) := (wbPartMux(197) xor i_prn(98)) & (not wbPartMux(196) xor i_prn(98)) & '1';
    wbMult(299 downto 297) := (wbPartMux(199) xor i_prn(99)) & (not wbPartMux(198) xor i_prn(99)) & '1';
    wbMult(302 downto 300) := (wbPartMux(201) xor i_prn(100)) & (not wbPartMux(200) xor i_prn(100)) & '1';
    wbMult(305 downto 303) := (wbPartMux(203) xor i_prn(101)) & (not wbPartMux(202) xor i_prn(101)) & '1';
    wbMult(308 downto 306) := (wbPartMux(205) xor i_prn(102)) & (not wbPartMux(204) xor i_prn(102)) & '1';
    wbMult(311 downto 309) := (wbPartMux(207) xor i_prn(103)) & (not wbPartMux(206) xor i_prn(103)) & '1';
    wbMult(314 downto 312) := (wbPartMux(209) xor i_prn(104)) & (not wbPartMux(208) xor i_prn(104)) & '1';
    wbMult(317 downto 315) := (wbPartMux(211) xor i_prn(105)) & (not wbPartMux(210) xor i_prn(105)) & '1';
    wbMult(320 downto 318) := (wbPartMux(213) xor i_prn(106)) & (not wbPartMux(212) xor i_prn(106)) & '1';
    wbMult(323 downto 321) := (wbPartMux(215) xor i_prn(107)) & (not wbPartMux(214) xor i_prn(107)) & '1';
    wbMult(326 downto 324) := (wbPartMux(217) xor i_prn(108)) & (not wbPartMux(216) xor i_prn(108)) & '1';
    wbMult(329 downto 327) := (wbPartMux(219) xor i_prn(109)) & (not wbPartMux(218) xor i_prn(109)) & '1';
    wbMult(332 downto 330) := (wbPartMux(221) xor i_prn(110)) & (not wbPartMux(220) xor i_prn(110)) & '1';
    wbMult(335 downto 333) := (wbPartMux(223) xor i_prn(111)) & (not wbPartMux(222) xor i_prn(111)) & '1';
    wbMult(338 downto 336) := (wbPartMux(225) xor i_prn(112)) & (not wbPartMux(224) xor i_prn(112)) & '1';
    wbMult(341 downto 339) := (wbPartMux(227) xor i_prn(113)) & (not wbPartMux(226) xor i_prn(113)) & '1';
    wbMult(344 downto 342) := (wbPartMux(229) xor i_prn(114)) & (not wbPartMux(228) xor i_prn(114)) & '1';
    wbMult(347 downto 345) := (wbPartMux(231) xor i_prn(115)) & (not wbPartMux(230) xor i_prn(115)) & '1';
    wbMult(350 downto 348) := (wbPartMux(233) xor i_prn(116)) & (not wbPartMux(232) xor i_prn(116)) & '1';
    wbMult(353 downto 351) := (wbPartMux(235) xor i_prn(117)) & (not wbPartMux(234) xor i_prn(117)) & '1';
    wbMult(356 downto 354) := (wbPartMux(237) xor i_prn(118)) & (not wbPartMux(236) xor i_prn(118)) & '1';
    wbMult(359 downto 357) := (wbPartMux(239) xor i_prn(119)) & (not wbPartMux(238) xor i_prn(119)) & '1';
    wbMult(362 downto 360) := (wbPartMux(241) xor i_prn(120)) & (not wbPartMux(240) xor i_prn(120)) & '1';
    wbMult(365 downto 363) := (wbPartMux(243) xor i_prn(121)) & (not wbPartMux(242) xor i_prn(121)) & '1';
    wbMult(368 downto 366) := (wbPartMux(245) xor i_prn(122)) & (not wbPartMux(244) xor i_prn(122)) & '1';
    wbMult(371 downto 369) := (wbPartMux(247) xor i_prn(123)) & (not wbPartMux(246) xor i_prn(123)) & '1';
    wbMult(374 downto 372) := (wbPartMux(249) xor i_prn(124)) & (not wbPartMux(248) xor i_prn(124)) & '1';
    wbMult(377 downto 375) := (wbPartMux(251) xor i_prn(125)) & (not wbPartMux(250) xor i_prn(125)) & '1';
    wbMult(380 downto 378) := (wbPartMux(253) xor i_prn(126)) & (not wbPartMux(252) xor i_prn(126)) & '1';
    wbMult(383 downto 381) := (wbPartMux(255) xor i_prn(127)) & (not wbPartMux(254) xor i_prn(127)) & '1';
    wbMult(386 downto 384) := (wbPartMux(257) xor i_prn(128)) & (not wbPartMux(256) xor i_prn(128)) & '1';
    wbMult(389 downto 387) := (wbPartMux(259) xor i_prn(129)) & (not wbPartMux(258) xor i_prn(129)) & '1';
    wbMult(392 downto 390) := (wbPartMux(261) xor i_prn(130)) & (not wbPartMux(260) xor i_prn(130)) & '1';
    wbMult(395 downto 393) := (wbPartMux(263) xor i_prn(131)) & (not wbPartMux(262) xor i_prn(131)) & '1';
    wbMult(398 downto 396) := (wbPartMux(265) xor i_prn(132)) & (not wbPartMux(264) xor i_prn(132)) & '1';
    wbMult(401 downto 399) := (wbPartMux(267) xor i_prn(133)) & (not wbPartMux(266) xor i_prn(133)) & '1';
    wbMult(404 downto 402) := (wbPartMux(269) xor i_prn(134)) & (not wbPartMux(268) xor i_prn(134)) & '1';
    wbMult(407 downto 405) := (wbPartMux(271) xor i_prn(135)) & (not wbPartMux(270) xor i_prn(135)) & '1';
    wbMult(410 downto 408) := (wbPartMux(273) xor i_prn(136)) & (not wbPartMux(272) xor i_prn(136)) & '1';
    wbMult(413 downto 411) := (wbPartMux(275) xor i_prn(137)) & (not wbPartMux(274) xor i_prn(137)) & '1';
    wbMult(416 downto 414) := (wbPartMux(277) xor i_prn(138)) & (not wbPartMux(276) xor i_prn(138)) & '1';
    wbMult(419 downto 417) := (wbPartMux(279) xor i_prn(139)) & (not wbPartMux(278) xor i_prn(139)) & '1';
    wbMult(422 downto 420) := (wbPartMux(281) xor i_prn(140)) & (not wbPartMux(280) xor i_prn(140)) & '1';
    wbMult(425 downto 423) := (wbPartMux(283) xor i_prn(141)) & (not wbPartMux(282) xor i_prn(141)) & '1';
    wbMult(428 downto 426) := (wbPartMux(285) xor i_prn(142)) & (not wbPartMux(284) xor i_prn(142)) & '1';
    wbMult(431 downto 429) := (wbPartMux(287) xor i_prn(143)) & (not wbPartMux(286) xor i_prn(143)) & '1';
    wbMult(434 downto 432) := (wbPartMux(289) xor i_prn(144)) & (not wbPartMux(288) xor i_prn(144)) & '1';
    wbMult(437 downto 435) := (wbPartMux(291) xor i_prn(145)) & (not wbPartMux(290) xor i_prn(145)) & '1';
    wbMult(440 downto 438) := (wbPartMux(293) xor i_prn(146)) & (not wbPartMux(292) xor i_prn(146)) & '1';
    wbMult(443 downto 441) := (wbPartMux(295) xor i_prn(147)) & (not wbPartMux(294) xor i_prn(147)) & '1';
    wbMult(446 downto 444) := (wbPartMux(297) xor i_prn(148)) & (not wbPartMux(296) xor i_prn(148)) & '1';
    wbMult(449 downto 447) := (wbPartMux(299) xor i_prn(149)) & (not wbPartMux(298) xor i_prn(149)) & '1';
    wbMult(452 downto 450) := (wbPartMux(301) xor i_prn(150)) & (not wbPartMux(300) xor i_prn(150)) & '1';
    wbMult(455 downto 453) := (wbPartMux(303) xor i_prn(151)) & (not wbPartMux(302) xor i_prn(151)) & '1';
    wbMult(458 downto 456) := (wbPartMux(305) xor i_prn(152)) & (not wbPartMux(304) xor i_prn(152)) & '1';
    wbMult(461 downto 459) := (wbPartMux(307) xor i_prn(153)) & (not wbPartMux(306) xor i_prn(153)) & '1';
    wbMult(464 downto 462) := (wbPartMux(309) xor i_prn(154)) & (not wbPartMux(308) xor i_prn(154)) & '1';
    wbMult(467 downto 465) := (wbPartMux(311) xor i_prn(155)) & (not wbPartMux(310) xor i_prn(155)) & '1';
    wbMult(470 downto 468) := (wbPartMux(313) xor i_prn(156)) & (not wbPartMux(312) xor i_prn(156)) & '1';
    wbMult(473 downto 471) := (wbPartMux(315) xor i_prn(157)) & (not wbPartMux(314) xor i_prn(157)) & '1';
    wbMult(476 downto 474) := (wbPartMux(317) xor i_prn(158)) & (not wbPartMux(316) xor i_prn(158)) & '1';
    wbMult(479 downto 477) := (wbPartMux(319) xor i_prn(159)) & (not wbPartMux(318) xor i_prn(159)) & '1';
    wbMult(482 downto 480) := (wbPartMux(321) xor i_prn(160)) & (not wbPartMux(320) xor i_prn(160)) & '1';
    wbMult(485 downto 483) := (wbPartMux(323) xor i_prn(161)) & (not wbPartMux(322) xor i_prn(161)) & '1';
    wbMult(488 downto 486) := (wbPartMux(325) xor i_prn(162)) & (not wbPartMux(324) xor i_prn(162)) & '1';
    wbMult(491 downto 489) := (wbPartMux(327) xor i_prn(163)) & (not wbPartMux(326) xor i_prn(163)) & '1';
    wbMult(494 downto 492) := (wbPartMux(329) xor i_prn(164)) & (not wbPartMux(328) xor i_prn(164)) & '1';
    wbMult(497 downto 495) := (wbPartMux(331) xor i_prn(165)) & (not wbPartMux(330) xor i_prn(165)) & '1';
    wbMult(500 downto 498) := (wbPartMux(333) xor i_prn(166)) & (not wbPartMux(332) xor i_prn(166)) & '1';
    wbMult(503 downto 501) := (wbPartMux(335) xor i_prn(167)) & (not wbPartMux(334) xor i_prn(167)) & '1';
    wbMult(506 downto 504) := (wbPartMux(337) xor i_prn(168)) & (not wbPartMux(336) xor i_prn(168)) & '1';
    wbMult(509 downto 507) := (wbPartMux(339) xor i_prn(169)) & (not wbPartMux(338) xor i_prn(169)) & '1';
    wbMult(512 downto 510) := (wbPartMux(341) xor i_prn(170)) & (not wbPartMux(340) xor i_prn(170)) & '1';
    wbMult(515 downto 513) := (wbPartMux(343) xor i_prn(171)) & (not wbPartMux(342) xor i_prn(171)) & '1';
    wbMult(518 downto 516) := (wbPartMux(345) xor i_prn(172)) & (not wbPartMux(344) xor i_prn(172)) & '1';
    wbMult(521 downto 519) := (wbPartMux(347) xor i_prn(173)) & (not wbPartMux(346) xor i_prn(173)) & '1';
    wbMult(524 downto 522) := (wbPartMux(349) xor i_prn(174)) & (not wbPartMux(348) xor i_prn(174)) & '1';
    wbMult(527 downto 525) := (wbPartMux(351) xor i_prn(175)) & (not wbPartMux(350) xor i_prn(175)) & '1';
    wbMult(530 downto 528) := (wbPartMux(353) xor i_prn(176)) & (not wbPartMux(352) xor i_prn(176)) & '1';
    wbMult(533 downto 531) := (wbPartMux(355) xor i_prn(177)) & (not wbPartMux(354) xor i_prn(177)) & '1';
    wbMult(536 downto 534) := (wbPartMux(357) xor i_prn(178)) & (not wbPartMux(356) xor i_prn(178)) & '1';
    wbMult(539 downto 537) := (wbPartMux(359) xor i_prn(179)) & (not wbPartMux(358) xor i_prn(179)) & '1';
    wbMult(542 downto 540) := (wbPartMux(361) xor i_prn(180)) & (not wbPartMux(360) xor i_prn(180)) & '1';
    wbMult(545 downto 543) := (wbPartMux(363) xor i_prn(181)) & (not wbPartMux(362) xor i_prn(181)) & '1';
    wbMult(548 downto 546) := (wbPartMux(365) xor i_prn(182)) & (not wbPartMux(364) xor i_prn(182)) & '1';
    wbMult(551 downto 549) := (wbPartMux(367) xor i_prn(183)) & (not wbPartMux(366) xor i_prn(183)) & '1';
    wbMult(554 downto 552) := (wbPartMux(369) xor i_prn(184)) & (not wbPartMux(368) xor i_prn(184)) & '1';
    wbMult(557 downto 555) := (wbPartMux(371) xor i_prn(185)) & (not wbPartMux(370) xor i_prn(185)) & '1';
    wbMult(560 downto 558) := (wbPartMux(373) xor i_prn(186)) & (not wbPartMux(372) xor i_prn(186)) & '1';
    wbMult(563 downto 561) := (wbPartMux(375) xor i_prn(187)) & (not wbPartMux(374) xor i_prn(187)) & '1';
    wbMult(566 downto 564) := (wbPartMux(377) xor i_prn(188)) & (not wbPartMux(376) xor i_prn(188)) & '1';
    wbMult(569 downto 567) := (wbPartMux(379) xor i_prn(189)) & (not wbPartMux(378) xor i_prn(189)) & '1';
    wbMult(572 downto 570) := (wbPartMux(381) xor i_prn(190)) & (not wbPartMux(380) xor i_prn(190)) & '1';
    wbMult(575 downto 573) := (wbPartMux(383) xor i_prn(191)) & (not wbPartMux(382) xor i_prn(191)) & '1';
    wbMult(578 downto 576) := (wbPartMux(385) xor i_prn(192)) & (not wbPartMux(384) xor i_prn(192)) & '1';
    wbMult(581 downto 579) := (wbPartMux(387) xor i_prn(193)) & (not wbPartMux(386) xor i_prn(193)) & '1';
    wbMult(584 downto 582) := (wbPartMux(389) xor i_prn(194)) & (not wbPartMux(388) xor i_prn(194)) & '1';
    wbMult(587 downto 585) := (wbPartMux(391) xor i_prn(195)) & (not wbPartMux(390) xor i_prn(195)) & '1';
    wbMult(590 downto 588) := (wbPartMux(393) xor i_prn(196)) & (not wbPartMux(392) xor i_prn(196)) & '1';
    wbMult(593 downto 591) := (wbPartMux(395) xor i_prn(197)) & (not wbPartMux(394) xor i_prn(197)) & '1';
    wbMult(596 downto 594) := (wbPartMux(397) xor i_prn(198)) & (not wbPartMux(396) xor i_prn(198)) & '1';
    wbMult(599 downto 597) := (wbPartMux(399) xor i_prn(199)) & (not wbPartMux(398) xor i_prn(199)) & '1';
    wbMult(602 downto 600) := (wbPartMux(401) xor i_prn(200)) & (not wbPartMux(400) xor i_prn(200)) & '1';
    wbMult(605 downto 603) := (wbPartMux(403) xor i_prn(201)) & (not wbPartMux(402) xor i_prn(201)) & '1';
    wbMult(608 downto 606) := (wbPartMux(405) xor i_prn(202)) & (not wbPartMux(404) xor i_prn(202)) & '1';
    wbMult(611 downto 609) := (wbPartMux(407) xor i_prn(203)) & (not wbPartMux(406) xor i_prn(203)) & '1';
    wbMult(614 downto 612) := (wbPartMux(409) xor i_prn(204)) & (not wbPartMux(408) xor i_prn(204)) & '1';
    wbMult(617 downto 615) := (wbPartMux(411) xor i_prn(205)) & (not wbPartMux(410) xor i_prn(205)) & '1';
    wbMult(620 downto 618) := (wbPartMux(413) xor i_prn(206)) & (not wbPartMux(412) xor i_prn(206)) & '1';
    wbMult(623 downto 621) := (wbPartMux(415) xor i_prn(207)) & (not wbPartMux(414) xor i_prn(207)) & '1';
    wbMult(626 downto 624) := (wbPartMux(417) xor i_prn(208)) & (not wbPartMux(416) xor i_prn(208)) & '1';
    wbMult(629 downto 627) := (wbPartMux(419) xor i_prn(209)) & (not wbPartMux(418) xor i_prn(209)) & '1';
    wbMult(632 downto 630) := (wbPartMux(421) xor i_prn(210)) & (not wbPartMux(420) xor i_prn(210)) & '1';
    wbMult(635 downto 633) := (wbPartMux(423) xor i_prn(211)) & (not wbPartMux(422) xor i_prn(211)) & '1';
    wbMult(638 downto 636) := (wbPartMux(425) xor i_prn(212)) & (not wbPartMux(424) xor i_prn(212)) & '1';
    wbMult(641 downto 639) := (wbPartMux(427) xor i_prn(213)) & (not wbPartMux(426) xor i_prn(213)) & '1';
    wbMult(644 downto 642) := (wbPartMux(429) xor i_prn(214)) & (not wbPartMux(428) xor i_prn(214)) & '1';
    wbMult(647 downto 645) := (wbPartMux(431) xor i_prn(215)) & (not wbPartMux(430) xor i_prn(215)) & '1';
    wbMult(650 downto 648) := (wbPartMux(433) xor i_prn(216)) & (not wbPartMux(432) xor i_prn(216)) & '1';
    wbMult(653 downto 651) := (wbPartMux(435) xor i_prn(217)) & (not wbPartMux(434) xor i_prn(217)) & '1';
    wbMult(656 downto 654) := (wbPartMux(437) xor i_prn(218)) & (not wbPartMux(436) xor i_prn(218)) & '1';
    wbMult(659 downto 657) := (wbPartMux(439) xor i_prn(219)) & (not wbPartMux(438) xor i_prn(219)) & '1';
    wbMult(662 downto 660) := (wbPartMux(441) xor i_prn(220)) & (not wbPartMux(440) xor i_prn(220)) & '1';
    wbMult(665 downto 663) := (wbPartMux(443) xor i_prn(221)) & (not wbPartMux(442) xor i_prn(221)) & '1';
    wbMult(668 downto 666) := (wbPartMux(445) xor i_prn(222)) & (not wbPartMux(444) xor i_prn(222)) & '1';
    wbMult(671 downto 669) := (wbPartMux(447) xor i_prn(223)) & (not wbPartMux(446) xor i_prn(223)) & '1';
    wbMult(674 downto 672) := (wbPartMux(449) xor i_prn(224)) & (not wbPartMux(448) xor i_prn(224)) & '1';
    wbMult(677 downto 675) := (wbPartMux(451) xor i_prn(225)) & (not wbPartMux(450) xor i_prn(225)) & '1';
    wbMult(680 downto 678) := (wbPartMux(453) xor i_prn(226)) & (not wbPartMux(452) xor i_prn(226)) & '1';
    wbMult(683 downto 681) := (wbPartMux(455) xor i_prn(227)) & (not wbPartMux(454) xor i_prn(227)) & '1';
    wbMult(686 downto 684) := (wbPartMux(457) xor i_prn(228)) & (not wbPartMux(456) xor i_prn(228)) & '1';
    wbMult(689 downto 687) := (wbPartMux(459) xor i_prn(229)) & (not wbPartMux(458) xor i_prn(229)) & '1';
    wbMult(692 downto 690) := (wbPartMux(461) xor i_prn(230)) & (not wbPartMux(460) xor i_prn(230)) & '1';
    wbMult(695 downto 693) := (wbPartMux(463) xor i_prn(231)) & (not wbPartMux(462) xor i_prn(231)) & '1';
    wbMult(698 downto 696) := (wbPartMux(465) xor i_prn(232)) & (not wbPartMux(464) xor i_prn(232)) & '1';
    wbMult(701 downto 699) := (wbPartMux(467) xor i_prn(233)) & (not wbPartMux(466) xor i_prn(233)) & '1';
    wbMult(704 downto 702) := (wbPartMux(469) xor i_prn(234)) & (not wbPartMux(468) xor i_prn(234)) & '1';
    wbMult(707 downto 705) := (wbPartMux(471) xor i_prn(235)) & (not wbPartMux(470) xor i_prn(235)) & '1';
    wbMult(710 downto 708) := (wbPartMux(473) xor i_prn(236)) & (not wbPartMux(472) xor i_prn(236)) & '1';
    wbMult(713 downto 711) := (wbPartMux(475) xor i_prn(237)) & (not wbPartMux(474) xor i_prn(237)) & '1';
    wbMult(716 downto 714) := (wbPartMux(477) xor i_prn(238)) & (not wbPartMux(476) xor i_prn(238)) & '1';
    wbMult(719 downto 717) := (wbPartMux(479) xor i_prn(239)) & (not wbPartMux(478) xor i_prn(239)) & '1';
    wbMult(722 downto 720) := (wbPartMux(481) xor i_prn(240)) & (not wbPartMux(480) xor i_prn(240)) & '1';
    wbMult(725 downto 723) := (wbPartMux(483) xor i_prn(241)) & (not wbPartMux(482) xor i_prn(241)) & '1';
    wbMult(728 downto 726) := (wbPartMux(485) xor i_prn(242)) & (not wbPartMux(484) xor i_prn(242)) & '1';
    wbMult(731 downto 729) := (wbPartMux(487) xor i_prn(243)) & (not wbPartMux(486) xor i_prn(243)) & '1';
    wbMult(734 downto 732) := (wbPartMux(489) xor i_prn(244)) & (not wbPartMux(488) xor i_prn(244)) & '1';
    wbMult(737 downto 735) := (wbPartMux(491) xor i_prn(245)) & (not wbPartMux(490) xor i_prn(245)) & '1';
    wbMult(740 downto 738) := (wbPartMux(493) xor i_prn(246)) & (not wbPartMux(492) xor i_prn(246)) & '1';
    wbMult(743 downto 741) := (wbPartMux(495) xor i_prn(247)) & (not wbPartMux(494) xor i_prn(247)) & '1';
    wbMult(746 downto 744) := (wbPartMux(497) xor i_prn(248)) & (not wbPartMux(496) xor i_prn(248)) & '1';
    wbMult(749 downto 747) := (wbPartMux(499) xor i_prn(249)) & (not wbPartMux(498) xor i_prn(249)) & '1';
    wbMult(752 downto 750) := (wbPartMux(501) xor i_prn(250)) & (not wbPartMux(500) xor i_prn(250)) & '1';
    wbMult(755 downto 753) := (wbPartMux(503) xor i_prn(251)) & (not wbPartMux(502) xor i_prn(251)) & '1';
    wbMult(758 downto 756) := (wbPartMux(505) xor i_prn(252)) & (not wbPartMux(504) xor i_prn(252)) & '1';
    wbMult(761 downto 759) := (wbPartMux(507) xor i_prn(253)) & (not wbPartMux(506) xor i_prn(253)) & '1';
    wbMult(764 downto 762) := (wbPartMux(509) xor i_prn(254)) & (not wbPartMux(508) xor i_prn(254)) & '1';
    wbMult(767 downto 765) := (wbPartMux(511) xor i_prn(255)) & (not wbPartMux(510) xor i_prn(255)) & '1';
    wbMult(770 downto 768) := (wbPartMux(513) xor i_prn(256)) & (not wbPartMux(512) xor i_prn(256)) & '1';
    wbMult(773 downto 771) := (wbPartMux(515) xor i_prn(257)) & (not wbPartMux(514) xor i_prn(257)) & '1';
    wbMult(776 downto 774) := (wbPartMux(517) xor i_prn(258)) & (not wbPartMux(516) xor i_prn(258)) & '1';
    wbMult(779 downto 777) := (wbPartMux(519) xor i_prn(259)) & (not wbPartMux(518) xor i_prn(259)) & '1';
    wbMult(782 downto 780) := (wbPartMux(521) xor i_prn(260)) & (not wbPartMux(520) xor i_prn(260)) & '1';
    wbMult(785 downto 783) := (wbPartMux(523) xor i_prn(261)) & (not wbPartMux(522) xor i_prn(261)) & '1';
    wbMult(788 downto 786) := (wbPartMux(525) xor i_prn(262)) & (not wbPartMux(524) xor i_prn(262)) & '1';
    wbMult(791 downto 789) := (wbPartMux(527) xor i_prn(263)) & (not wbPartMux(526) xor i_prn(263)) & '1';
    wbMult(794 downto 792) := (wbPartMux(529) xor i_prn(264)) & (not wbPartMux(528) xor i_prn(264)) & '1';
    wbMult(797 downto 795) := (wbPartMux(531) xor i_prn(265)) & (not wbPartMux(530) xor i_prn(265)) & '1';
    wbMult(800 downto 798) := (wbPartMux(533) xor i_prn(266)) & (not wbPartMux(532) xor i_prn(266)) & '1';
    wbMult(803 downto 801) := (wbPartMux(535) xor i_prn(267)) & (not wbPartMux(534) xor i_prn(267)) & '1';
    wbMult(806 downto 804) := (wbPartMux(537) xor i_prn(268)) & (not wbPartMux(536) xor i_prn(268)) & '1';
    wbMult(809 downto 807) := (wbPartMux(539) xor i_prn(269)) & (not wbPartMux(538) xor i_prn(269)) & '1';
    wbMult(812 downto 810) := (wbPartMux(541) xor i_prn(270)) & (not wbPartMux(540) xor i_prn(270)) & '1';
    wbMult(815 downto 813) := (wbPartMux(543) xor i_prn(271)) & (not wbPartMux(542) xor i_prn(271)) & '1';
    wbMult(818 downto 816) := (wbPartMux(545) xor i_prn(272)) & (not wbPartMux(544) xor i_prn(272)) & '1';
    wbMult(821 downto 819) := (wbPartMux(547) xor i_prn(273)) & (not wbPartMux(546) xor i_prn(273)) & '1';
    wbMult(824 downto 822) := (wbPartMux(549) xor i_prn(274)) & (not wbPartMux(548) xor i_prn(274)) & '1';
    wbMult(827 downto 825) := (wbPartMux(551) xor i_prn(275)) & (not wbPartMux(550) xor i_prn(275)) & '1';
    wbMult(830 downto 828) := (wbPartMux(553) xor i_prn(276)) & (not wbPartMux(552) xor i_prn(276)) & '1';
    wbMult(833 downto 831) := (wbPartMux(555) xor i_prn(277)) & (not wbPartMux(554) xor i_prn(277)) & '1';
    wbMult(836 downto 834) := (wbPartMux(557) xor i_prn(278)) & (not wbPartMux(556) xor i_prn(278)) & '1';
    wbMult(839 downto 837) := (wbPartMux(559) xor i_prn(279)) & (not wbPartMux(558) xor i_prn(279)) & '1';
    wbMult(842 downto 840) := (wbPartMux(561) xor i_prn(280)) & (not wbPartMux(560) xor i_prn(280)) & '1';
    wbMult(845 downto 843) := (wbPartMux(563) xor i_prn(281)) & (not wbPartMux(562) xor i_prn(281)) & '1';
    wbMult(848 downto 846) := (wbPartMux(565) xor i_prn(282)) & (not wbPartMux(564) xor i_prn(282)) & '1';
    wbMult(851 downto 849) := (wbPartMux(567) xor i_prn(283)) & (not wbPartMux(566) xor i_prn(283)) & '1';
    wbMult(854 downto 852) := (wbPartMux(569) xor i_prn(284)) & (not wbPartMux(568) xor i_prn(284)) & '1';
    wbMult(857 downto 855) := (wbPartMux(571) xor i_prn(285)) & (not wbPartMux(570) xor i_prn(285)) & '1';
    wbMult(860 downto 858) := (wbPartMux(573) xor i_prn(286)) & (not wbPartMux(572) xor i_prn(286)) & '1';
    wbMult(863 downto 861) := (wbPartMux(575) xor i_prn(287)) & (not wbPartMux(574) xor i_prn(287)) & '1';
    wbMult(866 downto 864) := (wbPartMux(577) xor i_prn(288)) & (not wbPartMux(576) xor i_prn(288)) & '1';
    wbMult(869 downto 867) := (wbPartMux(579) xor i_prn(289)) & (not wbPartMux(578) xor i_prn(289)) & '1';
    wbMult(872 downto 870) := (wbPartMux(581) xor i_prn(290)) & (not wbPartMux(580) xor i_prn(290)) & '1';
    wbMult(875 downto 873) := (wbPartMux(583) xor i_prn(291)) & (not wbPartMux(582) xor i_prn(291)) & '1';
    wbMult(878 downto 876) := (wbPartMux(585) xor i_prn(292)) & (not wbPartMux(584) xor i_prn(292)) & '1';
    wbMult(881 downto 879) := (wbPartMux(587) xor i_prn(293)) & (not wbPartMux(586) xor i_prn(293)) & '1';
    wbMult(884 downto 882) := (wbPartMux(589) xor i_prn(294)) & (not wbPartMux(588) xor i_prn(294)) & '1';
    wbMult(887 downto 885) := (wbPartMux(591) xor i_prn(295)) & (not wbPartMux(590) xor i_prn(295)) & '1';
    wbMult(890 downto 888) := (wbPartMux(593) xor i_prn(296)) & (not wbPartMux(592) xor i_prn(296)) & '1';
    wbMult(893 downto 891) := (wbPartMux(595) xor i_prn(297)) & (not wbPartMux(594) xor i_prn(297)) & '1';
    wbMult(896 downto 894) := (wbPartMux(597) xor i_prn(298)) & (not wbPartMux(596) xor i_prn(298)) & '1';
    wbMult(899 downto 897) := (wbPartMux(599) xor i_prn(299)) & (not wbPartMux(598) xor i_prn(299)) & '1';
    wbMult(902 downto 900) := (wbPartMux(601) xor i_prn(300)) & (not wbPartMux(600) xor i_prn(300)) & '1';
    wbMult(905 downto 903) := (wbPartMux(603) xor i_prn(301)) & (not wbPartMux(602) xor i_prn(301)) & '1';
    wbMult(908 downto 906) := (wbPartMux(605) xor i_prn(302)) & (not wbPartMux(604) xor i_prn(302)) & '1';
    wbMult(911 downto 909) := (wbPartMux(607) xor i_prn(303)) & (not wbPartMux(606) xor i_prn(303)) & '1';
    wbMult(914 downto 912) := (wbPartMux(609) xor i_prn(304)) & (not wbPartMux(608) xor i_prn(304)) & '1';
    wbMult(917 downto 915) := (wbPartMux(611) xor i_prn(305)) & (not wbPartMux(610) xor i_prn(305)) & '1';
    wbMult(920 downto 918) := (wbPartMux(613) xor i_prn(306)) & (not wbPartMux(612) xor i_prn(306)) & '1';
    wbMult(923 downto 921) := (wbPartMux(615) xor i_prn(307)) & (not wbPartMux(614) xor i_prn(307)) & '1';
    wbMult(926 downto 924) := (wbPartMux(617) xor i_prn(308)) & (not wbPartMux(616) xor i_prn(308)) & '1';
    wbMult(929 downto 927) := (wbPartMux(619) xor i_prn(309)) & (not wbPartMux(618) xor i_prn(309)) & '1';
    wbMult(932 downto 930) := (wbPartMux(621) xor i_prn(310)) & (not wbPartMux(620) xor i_prn(310)) & '1';
    wbMult(935 downto 933) := (wbPartMux(623) xor i_prn(311)) & (not wbPartMux(622) xor i_prn(311)) & '1';
    wbMult(938 downto 936) := (wbPartMux(625) xor i_prn(312)) & (not wbPartMux(624) xor i_prn(312)) & '1';
    wbMult(941 downto 939) := (wbPartMux(627) xor i_prn(313)) & (not wbPartMux(626) xor i_prn(313)) & '1';
    wbMult(944 downto 942) := (wbPartMux(629) xor i_prn(314)) & (not wbPartMux(628) xor i_prn(314)) & '1';
    wbMult(947 downto 945) := (wbPartMux(631) xor i_prn(315)) & (not wbPartMux(630) xor i_prn(315)) & '1';
    wbMult(950 downto 948) := (wbPartMux(633) xor i_prn(316)) & (not wbPartMux(632) xor i_prn(316)) & '1';
    wbMult(953 downto 951) := (wbPartMux(635) xor i_prn(317)) & (not wbPartMux(634) xor i_prn(317)) & '1';
    wbMult(956 downto 954) := (wbPartMux(637) xor i_prn(318)) & (not wbPartMux(636) xor i_prn(318)) & '1';
    wbMult(959 downto 957) := (wbPartMux(639) xor i_prn(319)) & (not wbPartMux(638) xor i_prn(319)) & '1';
    wbMult(962 downto 960) := (wbPartMux(641) xor i_prn(320)) & (not wbPartMux(640) xor i_prn(320)) & '1';
    wbMult(965 downto 963) := (wbPartMux(643) xor i_prn(321)) & (not wbPartMux(642) xor i_prn(321)) & '1';
    wbMult(968 downto 966) := (wbPartMux(645) xor i_prn(322)) & (not wbPartMux(644) xor i_prn(322)) & '1';
    wbMult(971 downto 969) := (wbPartMux(647) xor i_prn(323)) & (not wbPartMux(646) xor i_prn(323)) & '1';
    wbMult(974 downto 972) := (wbPartMux(649) xor i_prn(324)) & (not wbPartMux(648) xor i_prn(324)) & '1';
    wbMult(977 downto 975) := (wbPartMux(651) xor i_prn(325)) & (not wbPartMux(650) xor i_prn(325)) & '1';
    wbMult(980 downto 978) := (wbPartMux(653) xor i_prn(326)) & (not wbPartMux(652) xor i_prn(326)) & '1';
    wbMult(983 downto 981) := (wbPartMux(655) xor i_prn(327)) & (not wbPartMux(654) xor i_prn(327)) & '1';
    wbMult(986 downto 984) := (wbPartMux(657) xor i_prn(328)) & (not wbPartMux(656) xor i_prn(328)) & '1';
    wbMult(989 downto 987) := (wbPartMux(659) xor i_prn(329)) & (not wbPartMux(658) xor i_prn(329)) & '1';
    wbMult(992 downto 990) := (wbPartMux(661) xor i_prn(330)) & (not wbPartMux(660) xor i_prn(330)) & '1';
    wbMult(995 downto 993) := (wbPartMux(663) xor i_prn(331)) & (not wbPartMux(662) xor i_prn(331)) & '1';
    wbMult(998 downto 996) := (wbPartMux(665) xor i_prn(332)) & (not wbPartMux(664) xor i_prn(332)) & '1';
    wbMult(1001 downto 999) := (wbPartMux(667) xor i_prn(333)) & (not wbPartMux(666) xor i_prn(333)) & '1';
    wbMult(1004 downto 1002) := (wbPartMux(669) xor i_prn(334)) & (not wbPartMux(668) xor i_prn(334)) & '1';
    wbMult(1007 downto 1005) := (wbPartMux(671) xor i_prn(335)) & (not wbPartMux(670) xor i_prn(335)) & '1';
    wbMult(1010 downto 1008) := (wbPartMux(673) xor i_prn(336)) & (not wbPartMux(672) xor i_prn(336)) & '1';
    wbMult(1013 downto 1011) := (wbPartMux(675) xor i_prn(337)) & (not wbPartMux(674) xor i_prn(337)) & '1';
    wbMult(1016 downto 1014) := (wbPartMux(677) xor i_prn(338)) & (not wbPartMux(676) xor i_prn(338)) & '1';
    wbMult(1019 downto 1017) := (wbPartMux(679) xor i_prn(339)) & (not wbPartMux(678) xor i_prn(339)) & '1';
    wbMult(1022 downto 1020) := (wbPartMux(681) xor i_prn(340)) & (not wbPartMux(680) xor i_prn(340)) & '1';
    wbMult(1025 downto 1023) := (wbPartMux(683) xor i_prn(341)) & (not wbPartMux(682) xor i_prn(341)) & '1';
    wbMult(1028 downto 1026) := (wbPartMux(685) xor i_prn(342)) & (not wbPartMux(684) xor i_prn(342)) & '1';
    wbMult(1031 downto 1029) := (wbPartMux(687) xor i_prn(343)) & (not wbPartMux(686) xor i_prn(343)) & '1';
    wbMult(1034 downto 1032) := (wbPartMux(689) xor i_prn(344)) & (not wbPartMux(688) xor i_prn(344)) & '1';
    wbMult(1037 downto 1035) := (wbPartMux(691) xor i_prn(345)) & (not wbPartMux(690) xor i_prn(345)) & '1';
    wbMult(1040 downto 1038) := (wbPartMux(693) xor i_prn(346)) & (not wbPartMux(692) xor i_prn(346)) & '1';
    wbMult(1043 downto 1041) := (wbPartMux(695) xor i_prn(347)) & (not wbPartMux(694) xor i_prn(347)) & '1';
    wbMult(1046 downto 1044) := (wbPartMux(697) xor i_prn(348)) & (not wbPartMux(696) xor i_prn(348)) & '1';
    wbMult(1049 downto 1047) := (wbPartMux(699) xor i_prn(349)) & (not wbPartMux(698) xor i_prn(349)) & '1';
    wbMult(1052 downto 1050) := (wbPartMux(701) xor i_prn(350)) & (not wbPartMux(700) xor i_prn(350)) & '1';
    wbMult(1055 downto 1053) := (wbPartMux(703) xor i_prn(351)) & (not wbPartMux(702) xor i_prn(351)) & '1';
    wbMult(1058 downto 1056) := (wbPartMux(705) xor i_prn(352)) & (not wbPartMux(704) xor i_prn(352)) & '1';
    wbMult(1061 downto 1059) := (wbPartMux(707) xor i_prn(353)) & (not wbPartMux(706) xor i_prn(353)) & '1';
    wbMult(1064 downto 1062) := (wbPartMux(709) xor i_prn(354)) & (not wbPartMux(708) xor i_prn(354)) & '1';
    wbMult(1067 downto 1065) := (wbPartMux(711) xor i_prn(355)) & (not wbPartMux(710) xor i_prn(355)) & '1';
    wbMult(1070 downto 1068) := (wbPartMux(713) xor i_prn(356)) & (not wbPartMux(712) xor i_prn(356)) & '1';
    wbMult(1073 downto 1071) := (wbPartMux(715) xor i_prn(357)) & (not wbPartMux(714) xor i_prn(357)) & '1';
    wbMult(1076 downto 1074) := (wbPartMux(717) xor i_prn(358)) & (not wbPartMux(716) xor i_prn(358)) & '1';
    wbMult(1079 downto 1077) := (wbPartMux(719) xor i_prn(359)) & (not wbPartMux(718) xor i_prn(359)) & '1';
    wbMult(1082 downto 1080) := (wbPartMux(721) xor i_prn(360)) & (not wbPartMux(720) xor i_prn(360)) & '1';
    wbMult(1085 downto 1083) := (wbPartMux(723) xor i_prn(361)) & (not wbPartMux(722) xor i_prn(361)) & '1';
    wbMult(1088 downto 1086) := (wbPartMux(725) xor i_prn(362)) & (not wbPartMux(724) xor i_prn(362)) & '1';
    wbMult(1091 downto 1089) := (wbPartMux(727) xor i_prn(363)) & (not wbPartMux(726) xor i_prn(363)) & '1';
    wbMult(1094 downto 1092) := (wbPartMux(729) xor i_prn(364)) & (not wbPartMux(728) xor i_prn(364)) & '1';
    wbMult(1097 downto 1095) := (wbPartMux(731) xor i_prn(365)) & (not wbPartMux(730) xor i_prn(365)) & '1';
    wbMult(1100 downto 1098) := (wbPartMux(733) xor i_prn(366)) & (not wbPartMux(732) xor i_prn(366)) & '1';
    wbMult(1103 downto 1101) := (wbPartMux(735) xor i_prn(367)) & (not wbPartMux(734) xor i_prn(367)) & '1';
    wbMult(1106 downto 1104) := (wbPartMux(737) xor i_prn(368)) & (not wbPartMux(736) xor i_prn(368)) & '1';
    wbMult(1109 downto 1107) := (wbPartMux(739) xor i_prn(369)) & (not wbPartMux(738) xor i_prn(369)) & '1';
    wbMult(1112 downto 1110) := (wbPartMux(741) xor i_prn(370)) & (not wbPartMux(740) xor i_prn(370)) & '1';
    wbMult(1115 downto 1113) := (wbPartMux(743) xor i_prn(371)) & (not wbPartMux(742) xor i_prn(371)) & '1';
    wbMult(1118 downto 1116) := (wbPartMux(745) xor i_prn(372)) & (not wbPartMux(744) xor i_prn(372)) & '1';
    wbMult(1121 downto 1119) := (wbPartMux(747) xor i_prn(373)) & (not wbPartMux(746) xor i_prn(373)) & '1';
    wbMult(1124 downto 1122) := (wbPartMux(749) xor i_prn(374)) & (not wbPartMux(748) xor i_prn(374)) & '1';
    wbMult(1127 downto 1125) := (wbPartMux(751) xor i_prn(375)) & (not wbPartMux(750) xor i_prn(375)) & '1';
    wbMult(1130 downto 1128) := (wbPartMux(753) xor i_prn(376)) & (not wbPartMux(752) xor i_prn(376)) & '1';
    wbMult(1133 downto 1131) := (wbPartMux(755) xor i_prn(377)) & (not wbPartMux(754) xor i_prn(377)) & '1';
    wbMult(1136 downto 1134) := (wbPartMux(757) xor i_prn(378)) & (not wbPartMux(756) xor i_prn(378)) & '1';
    wbMult(1139 downto 1137) := (wbPartMux(759) xor i_prn(379)) & (not wbPartMux(758) xor i_prn(379)) & '1';
    wbMult(1142 downto 1140) := (wbPartMux(761) xor i_prn(380)) & (not wbPartMux(760) xor i_prn(380)) & '1';
    wbMult(1145 downto 1143) := (wbPartMux(763) xor i_prn(381)) & (not wbPartMux(762) xor i_prn(381)) & '1';
    wbMult(1148 downto 1146) := (wbPartMux(765) xor i_prn(382)) & (not wbPartMux(764) xor i_prn(382)) & '1';
    wbMult(1151 downto 1149) := (wbPartMux(767) xor i_prn(383)) & (not wbPartMux(766) xor i_prn(383)) & '1';
    wbMult(1154 downto 1152) := (wbPartMux(769) xor i_prn(384)) & (not wbPartMux(768) xor i_prn(384)) & '1';
    wbMult(1157 downto 1155) := (wbPartMux(771) xor i_prn(385)) & (not wbPartMux(770) xor i_prn(385)) & '1';
    wbMult(1160 downto 1158) := (wbPartMux(773) xor i_prn(386)) & (not wbPartMux(772) xor i_prn(386)) & '1';
    wbMult(1163 downto 1161) := (wbPartMux(775) xor i_prn(387)) & (not wbPartMux(774) xor i_prn(387)) & '1';
    wbMult(1166 downto 1164) := (wbPartMux(777) xor i_prn(388)) & (not wbPartMux(776) xor i_prn(388)) & '1';
    wbMult(1169 downto 1167) := (wbPartMux(779) xor i_prn(389)) & (not wbPartMux(778) xor i_prn(389)) & '1';
    wbMult(1172 downto 1170) := (wbPartMux(781) xor i_prn(390)) & (not wbPartMux(780) xor i_prn(390)) & '1';
    wbMult(1175 downto 1173) := (wbPartMux(783) xor i_prn(391)) & (not wbPartMux(782) xor i_prn(391)) & '1';
    wbMult(1178 downto 1176) := (wbPartMux(785) xor i_prn(392)) & (not wbPartMux(784) xor i_prn(392)) & '1';
    wbMult(1181 downto 1179) := (wbPartMux(787) xor i_prn(393)) & (not wbPartMux(786) xor i_prn(393)) & '1';
    wbMult(1184 downto 1182) := (wbPartMux(789) xor i_prn(394)) & (not wbPartMux(788) xor i_prn(394)) & '1';
    wbMult(1187 downto 1185) := (wbPartMux(791) xor i_prn(395)) & (not wbPartMux(790) xor i_prn(395)) & '1';
    wbMult(1190 downto 1188) := (wbPartMux(793) xor i_prn(396)) & (not wbPartMux(792) xor i_prn(396)) & '1';
    wbMult(1193 downto 1191) := (wbPartMux(795) xor i_prn(397)) & (not wbPartMux(794) xor i_prn(397)) & '1';
    wbMult(1196 downto 1194) := (wbPartMux(797) xor i_prn(398)) & (not wbPartMux(796) xor i_prn(398)) & '1';
    wbMult(1199 downto 1197) := (wbPartMux(799) xor i_prn(399)) & (not wbPartMux(798) xor i_prn(399)) & '1';
    wbMult(1202 downto 1200) := (wbPartMux(801) xor i_prn(400)) & (not wbPartMux(800) xor i_prn(400)) & '1';
    wbMult(1205 downto 1203) := (wbPartMux(803) xor i_prn(401)) & (not wbPartMux(802) xor i_prn(401)) & '1';
    wbMult(1208 downto 1206) := (wbPartMux(805) xor i_prn(402)) & (not wbPartMux(804) xor i_prn(402)) & '1';
    wbMult(1211 downto 1209) := (wbPartMux(807) xor i_prn(403)) & (not wbPartMux(806) xor i_prn(403)) & '1';
    wbMult(1214 downto 1212) := (wbPartMux(809) xor i_prn(404)) & (not wbPartMux(808) xor i_prn(404)) & '1';
    wbMult(1217 downto 1215) := (wbPartMux(811) xor i_prn(405)) & (not wbPartMux(810) xor i_prn(405)) & '1';
    wbMult(1220 downto 1218) := (wbPartMux(813) xor i_prn(406)) & (not wbPartMux(812) xor i_prn(406)) & '1';
    wbMult(1223 downto 1221) := (wbPartMux(815) xor i_prn(407)) & (not wbPartMux(814) xor i_prn(407)) & '1';
    wbMult(1226 downto 1224) := (wbPartMux(817) xor i_prn(408)) & (not wbPartMux(816) xor i_prn(408)) & '1';
    wbMult(1229 downto 1227) := (wbPartMux(819) xor i_prn(409)) & (not wbPartMux(818) xor i_prn(409)) & '1';
    wbMult(1232 downto 1230) := (wbPartMux(821) xor i_prn(410)) & (not wbPartMux(820) xor i_prn(410)) & '1';
    wbMult(1235 downto 1233) := (wbPartMux(823) xor i_prn(411)) & (not wbPartMux(822) xor i_prn(411)) & '1';
    wbMult(1238 downto 1236) := (wbPartMux(825) xor i_prn(412)) & (not wbPartMux(824) xor i_prn(412)) & '1';
    wbMult(1241 downto 1239) := (wbPartMux(827) xor i_prn(413)) & (not wbPartMux(826) xor i_prn(413)) & '1';
    wbMult(1244 downto 1242) := (wbPartMux(829) xor i_prn(414)) & (not wbPartMux(828) xor i_prn(414)) & '1';
    wbMult(1247 downto 1245) := (wbPartMux(831) xor i_prn(415)) & (not wbPartMux(830) xor i_prn(415)) & '1';
    wbMult(1250 downto 1248) := (wbPartMux(833) xor i_prn(416)) & (not wbPartMux(832) xor i_prn(416)) & '1';
    wbMult(1253 downto 1251) := (wbPartMux(835) xor i_prn(417)) & (not wbPartMux(834) xor i_prn(417)) & '1';
    wbMult(1256 downto 1254) := (wbPartMux(837) xor i_prn(418)) & (not wbPartMux(836) xor i_prn(418)) & '1';
    wbMult(1259 downto 1257) := (wbPartMux(839) xor i_prn(419)) & (not wbPartMux(838) xor i_prn(419)) & '1';
    wbMult(1262 downto 1260) := (wbPartMux(841) xor i_prn(420)) & (not wbPartMux(840) xor i_prn(420)) & '1';
    wbMult(1265 downto 1263) := (wbPartMux(843) xor i_prn(421)) & (not wbPartMux(842) xor i_prn(421)) & '1';
    wbMult(1268 downto 1266) := (wbPartMux(845) xor i_prn(422)) & (not wbPartMux(844) xor i_prn(422)) & '1';
    wbMult(1271 downto 1269) := (wbPartMux(847) xor i_prn(423)) & (not wbPartMux(846) xor i_prn(423)) & '1';
    wbMult(1274 downto 1272) := (wbPartMux(849) xor i_prn(424)) & (not wbPartMux(848) xor i_prn(424)) & '1';
    wbMult(1277 downto 1275) := (wbPartMux(851) xor i_prn(425)) & (not wbPartMux(850) xor i_prn(425)) & '1';
    wbMult(1280 downto 1278) := (wbPartMux(853) xor i_prn(426)) & (not wbPartMux(852) xor i_prn(426)) & '1';
    wbMult(1283 downto 1281) := (wbPartMux(855) xor i_prn(427)) & (not wbPartMux(854) xor i_prn(427)) & '1';
    wbMult(1286 downto 1284) := (wbPartMux(857) xor i_prn(428)) & (not wbPartMux(856) xor i_prn(428)) & '1';
    wbMult(1289 downto 1287) := (wbPartMux(859) xor i_prn(429)) & (not wbPartMux(858) xor i_prn(429)) & '1';
    wbMult(1292 downto 1290) := (wbPartMux(861) xor i_prn(430)) & (not wbPartMux(860) xor i_prn(430)) & '1';
    wbMult(1295 downto 1293) := (wbPartMux(863) xor i_prn(431)) & (not wbPartMux(862) xor i_prn(431)) & '1';
    wbMult(1298 downto 1296) := (wbPartMux(865) xor i_prn(432)) & (not wbPartMux(864) xor i_prn(432)) & '1';
    wbMult(1301 downto 1299) := (wbPartMux(867) xor i_prn(433)) & (not wbPartMux(866) xor i_prn(433)) & '1';
    wbMult(1304 downto 1302) := (wbPartMux(869) xor i_prn(434)) & (not wbPartMux(868) xor i_prn(434)) & '1';
    wbMult(1307 downto 1305) := (wbPartMux(871) xor i_prn(435)) & (not wbPartMux(870) xor i_prn(435)) & '1';
    wbMult(1310 downto 1308) := (wbPartMux(873) xor i_prn(436)) & (not wbPartMux(872) xor i_prn(436)) & '1';
    wbMult(1313 downto 1311) := (wbPartMux(875) xor i_prn(437)) & (not wbPartMux(874) xor i_prn(437)) & '1';
    wbMult(1316 downto 1314) := (wbPartMux(877) xor i_prn(438)) & (not wbPartMux(876) xor i_prn(438)) & '1';
    wbMult(1319 downto 1317) := (wbPartMux(879) xor i_prn(439)) & (not wbPartMux(878) xor i_prn(439)) & '1';
    wbMult(1322 downto 1320) := (wbPartMux(881) xor i_prn(440)) & (not wbPartMux(880) xor i_prn(440)) & '1';
    wbMult(1325 downto 1323) := (wbPartMux(883) xor i_prn(441)) & (not wbPartMux(882) xor i_prn(441)) & '1';
    wbMult(1328 downto 1326) := (wbPartMux(885) xor i_prn(442)) & (not wbPartMux(884) xor i_prn(442)) & '1';
    wbMult(1331 downto 1329) := (wbPartMux(887) xor i_prn(443)) & (not wbPartMux(886) xor i_prn(443)) & '1';
    wbMult(1334 downto 1332) := (wbPartMux(889) xor i_prn(444)) & (not wbPartMux(888) xor i_prn(444)) & '1';
    wbMult(1337 downto 1335) := (wbPartMux(891) xor i_prn(445)) & (not wbPartMux(890) xor i_prn(445)) & '1';
    wbMult(1340 downto 1338) := (wbPartMux(893) xor i_prn(446)) & (not wbPartMux(892) xor i_prn(446)) & '1';
    wbMult(1343 downto 1341) := (wbPartMux(895) xor i_prn(447)) & (not wbPartMux(894) xor i_prn(447)) & '1';
    wbMult(1346 downto 1344) := (wbPartMux(897) xor i_prn(448)) & (not wbPartMux(896) xor i_prn(448)) & '1';
    wbMult(1349 downto 1347) := (wbPartMux(899) xor i_prn(449)) & (not wbPartMux(898) xor i_prn(449)) & '1';
    wbMult(1352 downto 1350) := (wbPartMux(901) xor i_prn(450)) & (not wbPartMux(900) xor i_prn(450)) & '1';
    wbMult(1355 downto 1353) := (wbPartMux(903) xor i_prn(451)) & (not wbPartMux(902) xor i_prn(451)) & '1';
    wbMult(1358 downto 1356) := (wbPartMux(905) xor i_prn(452)) & (not wbPartMux(904) xor i_prn(452)) & '1';
    wbMult(1361 downto 1359) := (wbPartMux(907) xor i_prn(453)) & (not wbPartMux(906) xor i_prn(453)) & '1';
    wbMult(1364 downto 1362) := (wbPartMux(909) xor i_prn(454)) & (not wbPartMux(908) xor i_prn(454)) & '1';
    wbMult(1367 downto 1365) := (wbPartMux(911) xor i_prn(455)) & (not wbPartMux(910) xor i_prn(455)) & '1';
    wbMult(1370 downto 1368) := (wbPartMux(913) xor i_prn(456)) & (not wbPartMux(912) xor i_prn(456)) & '1';
    wbMult(1373 downto 1371) := (wbPartMux(915) xor i_prn(457)) & (not wbPartMux(914) xor i_prn(457)) & '1';
    wbMult(1376 downto 1374) := (wbPartMux(917) xor i_prn(458)) & (not wbPartMux(916) xor i_prn(458)) & '1';
    wbMult(1379 downto 1377) := (wbPartMux(919) xor i_prn(459)) & (not wbPartMux(918) xor i_prn(459)) & '1';
    wbMult(1382 downto 1380) := (wbPartMux(921) xor i_prn(460)) & (not wbPartMux(920) xor i_prn(460)) & '1';
    wbMult(1385 downto 1383) := (wbPartMux(923) xor i_prn(461)) & (not wbPartMux(922) xor i_prn(461)) & '1';
    wbMult(1388 downto 1386) := (wbPartMux(925) xor i_prn(462)) & (not wbPartMux(924) xor i_prn(462)) & '1';
    wbMult(1391 downto 1389) := (wbPartMux(927) xor i_prn(463)) & (not wbPartMux(926) xor i_prn(463)) & '1';
    wbMult(1394 downto 1392) := (wbPartMux(929) xor i_prn(464)) & (not wbPartMux(928) xor i_prn(464)) & '1';
    wbMult(1397 downto 1395) := (wbPartMux(931) xor i_prn(465)) & (not wbPartMux(930) xor i_prn(465)) & '1';
    wbMult(1400 downto 1398) := (wbPartMux(933) xor i_prn(466)) & (not wbPartMux(932) xor i_prn(466)) & '1';
    wbMult(1403 downto 1401) := (wbPartMux(935) xor i_prn(467)) & (not wbPartMux(934) xor i_prn(467)) & '1';
    wbMult(1406 downto 1404) := (wbPartMux(937) xor i_prn(468)) & (not wbPartMux(936) xor i_prn(468)) & '1';
    wbMult(1409 downto 1407) := (wbPartMux(939) xor i_prn(469)) & (not wbPartMux(938) xor i_prn(469)) & '1';
    wbMult(1412 downto 1410) := (wbPartMux(941) xor i_prn(470)) & (not wbPartMux(940) xor i_prn(470)) & '1';
    wbMult(1415 downto 1413) := (wbPartMux(943) xor i_prn(471)) & (not wbPartMux(942) xor i_prn(471)) & '1';
    wbMult(1418 downto 1416) := (wbPartMux(945) xor i_prn(472)) & (not wbPartMux(944) xor i_prn(472)) & '1';
    wbMult(1421 downto 1419) := (wbPartMux(947) xor i_prn(473)) & (not wbPartMux(946) xor i_prn(473)) & '1';
    wbMult(1424 downto 1422) := (wbPartMux(949) xor i_prn(474)) & (not wbPartMux(948) xor i_prn(474)) & '1';
    wbMult(1427 downto 1425) := (wbPartMux(951) xor i_prn(475)) & (not wbPartMux(950) xor i_prn(475)) & '1';
    wbMult(1430 downto 1428) := (wbPartMux(953) xor i_prn(476)) & (not wbPartMux(952) xor i_prn(476)) & '1';
    wbMult(1433 downto 1431) := (wbPartMux(955) xor i_prn(477)) & (not wbPartMux(954) xor i_prn(477)) & '1';
    wbMult(1436 downto 1434) := (wbPartMux(957) xor i_prn(478)) & (not wbPartMux(956) xor i_prn(478)) & '1';
    wbMult(1439 downto 1437) := (wbPartMux(959) xor i_prn(479)) & (not wbPartMux(958) xor i_prn(479)) & '1';
    wbMult(1442 downto 1440) := (wbPartMux(961) xor i_prn(480)) & (not wbPartMux(960) xor i_prn(480)) & '1';
    wbMult(1445 downto 1443) := (wbPartMux(963) xor i_prn(481)) & (not wbPartMux(962) xor i_prn(481)) & '1';
    wbMult(1448 downto 1446) := (wbPartMux(965) xor i_prn(482)) & (not wbPartMux(964) xor i_prn(482)) & '1';
    wbMult(1451 downto 1449) := (wbPartMux(967) xor i_prn(483)) & (not wbPartMux(966) xor i_prn(483)) & '1';
    wbMult(1454 downto 1452) := (wbPartMux(969) xor i_prn(484)) & (not wbPartMux(968) xor i_prn(484)) & '1';
    wbMult(1457 downto 1455) := (wbPartMux(971) xor i_prn(485)) & (not wbPartMux(970) xor i_prn(485)) & '1';
    wbMult(1460 downto 1458) := (wbPartMux(973) xor i_prn(486)) & (not wbPartMux(972) xor i_prn(486)) & '1';
    wbMult(1463 downto 1461) := (wbPartMux(975) xor i_prn(487)) & (not wbPartMux(974) xor i_prn(487)) & '1';
    wbMult(1466 downto 1464) := (wbPartMux(977) xor i_prn(488)) & (not wbPartMux(976) xor i_prn(488)) & '1';
    wbMult(1469 downto 1467) := (wbPartMux(979) xor i_prn(489)) & (not wbPartMux(978) xor i_prn(489)) & '1';
    wbMult(1472 downto 1470) := (wbPartMux(981) xor i_prn(490)) & (not wbPartMux(980) xor i_prn(490)) & '1';
    wbMult(1475 downto 1473) := (wbPartMux(983) xor i_prn(491)) & (not wbPartMux(982) xor i_prn(491)) & '1';
    wbMult(1478 downto 1476) := (wbPartMux(985) xor i_prn(492)) & (not wbPartMux(984) xor i_prn(492)) & '1';
    wbMult(1481 downto 1479) := (wbPartMux(987) xor i_prn(493)) & (not wbPartMux(986) xor i_prn(493)) & '1';
    wbMult(1484 downto 1482) := (wbPartMux(989) xor i_prn(494)) & (not wbPartMux(988) xor i_prn(494)) & '1';
    wbMult(1487 downto 1485) := (wbPartMux(991) xor i_prn(495)) & (not wbPartMux(990) xor i_prn(495)) & '1';
    wbMult(1490 downto 1488) := (wbPartMux(993) xor i_prn(496)) & (not wbPartMux(992) xor i_prn(496)) & '1';
    wbMult(1493 downto 1491) := (wbPartMux(995) xor i_prn(497)) & (not wbPartMux(994) xor i_prn(497)) & '1';
    wbMult(1496 downto 1494) := (wbPartMux(997) xor i_prn(498)) & (not wbPartMux(996) xor i_prn(498)) & '1';
    wbMult(1499 downto 1497) := (wbPartMux(999) xor i_prn(499)) & (not wbPartMux(998) xor i_prn(499)) & '1';
    wbMult(1502 downto 1500) := (wbPartMux(1001) xor i_prn(500)) & (not wbPartMux(1000) xor i_prn(500)) & '1';
    wbMult(1505 downto 1503) := (wbPartMux(1003) xor i_prn(501)) & (not wbPartMux(1002) xor i_prn(501)) & '1';
    wbMult(1508 downto 1506) := (wbPartMux(1005) xor i_prn(502)) & (not wbPartMux(1004) xor i_prn(502)) & '1';
    wbMult(1511 downto 1509) := (wbPartMux(1007) xor i_prn(503)) & (not wbPartMux(1006) xor i_prn(503)) & '1';
    wbMult(1514 downto 1512) := (wbPartMux(1009) xor i_prn(504)) & (not wbPartMux(1008) xor i_prn(504)) & '1';
    wbMult(1517 downto 1515) := (wbPartMux(1011) xor i_prn(505)) & (not wbPartMux(1010) xor i_prn(505)) & '1';
    wbMult(1520 downto 1518) := (wbPartMux(1013) xor i_prn(506)) & (not wbPartMux(1012) xor i_prn(506)) & '1';
    wbMult(1523 downto 1521) := (wbPartMux(1015) xor i_prn(507)) & (not wbPartMux(1014) xor i_prn(507)) & '1';
    wbMult(1526 downto 1524) := (wbPartMux(1017) xor i_prn(508)) & (not wbPartMux(1016) xor i_prn(508)) & '1';
    wbMult(1529 downto 1527) := (wbPartMux(1019) xor i_prn(509)) & (not wbPartMux(1018) xor i_prn(509)) & '1';
    wbMult(1532 downto 1530) := (wbPartMux(1021) xor i_prn(510)) & (not wbPartMux(1020) xor i_prn(510)) & '1';
    wbMult(1535 downto 1533) := (wbPartMux(1023) xor i_prn(511)) & (not wbPartMux(1022) xor i_prn(511)) & '1';
    wbMult(1538 downto 1536) := (wbPartMux(1025) xor i_prn(512)) & (not wbPartMux(1024) xor i_prn(512)) & '1';
    wbMult(1541 downto 1539) := (wbPartMux(1027) xor i_prn(513)) & (not wbPartMux(1026) xor i_prn(513)) & '1';
    wbMult(1544 downto 1542) := (wbPartMux(1029) xor i_prn(514)) & (not wbPartMux(1028) xor i_prn(514)) & '1';
    wbMult(1547 downto 1545) := (wbPartMux(1031) xor i_prn(515)) & (not wbPartMux(1030) xor i_prn(515)) & '1';
    wbMult(1550 downto 1548) := (wbPartMux(1033) xor i_prn(516)) & (not wbPartMux(1032) xor i_prn(516)) & '1';
    wbMult(1553 downto 1551) := (wbPartMux(1035) xor i_prn(517)) & (not wbPartMux(1034) xor i_prn(517)) & '1';
    wbMult(1556 downto 1554) := (wbPartMux(1037) xor i_prn(518)) & (not wbPartMux(1036) xor i_prn(518)) & '1';
    wbMult(1559 downto 1557) := (wbPartMux(1039) xor i_prn(519)) & (not wbPartMux(1038) xor i_prn(519)) & '1';
    wbMult(1562 downto 1560) := (wbPartMux(1041) xor i_prn(520)) & (not wbPartMux(1040) xor i_prn(520)) & '1';
    wbMult(1565 downto 1563) := (wbPartMux(1043) xor i_prn(521)) & (not wbPartMux(1042) xor i_prn(521)) & '1';
    wbMult(1568 downto 1566) := (wbPartMux(1045) xor i_prn(522)) & (not wbPartMux(1044) xor i_prn(522)) & '1';
    wbMult(1571 downto 1569) := (wbPartMux(1047) xor i_prn(523)) & (not wbPartMux(1046) xor i_prn(523)) & '1';
    wbMult(1574 downto 1572) := (wbPartMux(1049) xor i_prn(524)) & (not wbPartMux(1048) xor i_prn(524)) & '1';
    wbMult(1577 downto 1575) := (wbPartMux(1051) xor i_prn(525)) & (not wbPartMux(1050) xor i_prn(525)) & '1';
    wbMult(1580 downto 1578) := (wbPartMux(1053) xor i_prn(526)) & (not wbPartMux(1052) xor i_prn(526)) & '1';
    wbMult(1583 downto 1581) := (wbPartMux(1055) xor i_prn(527)) & (not wbPartMux(1054) xor i_prn(527)) & '1';
    wbMult(1586 downto 1584) := (wbPartMux(1057) xor i_prn(528)) & (not wbPartMux(1056) xor i_prn(528)) & '1';
    wbMult(1589 downto 1587) := (wbPartMux(1059) xor i_prn(529)) & (not wbPartMux(1058) xor i_prn(529)) & '1';
    wbMult(1592 downto 1590) := (wbPartMux(1061) xor i_prn(530)) & (not wbPartMux(1060) xor i_prn(530)) & '1';
    wbMult(1595 downto 1593) := (wbPartMux(1063) xor i_prn(531)) & (not wbPartMux(1062) xor i_prn(531)) & '1';
    wbMult(1598 downto 1596) := (wbPartMux(1065) xor i_prn(532)) & (not wbPartMux(1064) xor i_prn(532)) & '1';
    wbMult(1601 downto 1599) := (wbPartMux(1067) xor i_prn(533)) & (not wbPartMux(1066) xor i_prn(533)) & '1';
    wbMult(1604 downto 1602) := (wbPartMux(1069) xor i_prn(534)) & (not wbPartMux(1068) xor i_prn(534)) & '1';
    wbMult(1607 downto 1605) := (wbPartMux(1071) xor i_prn(535)) & (not wbPartMux(1070) xor i_prn(535)) & '1';
    wbMult(1610 downto 1608) := (wbPartMux(1073) xor i_prn(536)) & (not wbPartMux(1072) xor i_prn(536)) & '1';
    wbMult(1613 downto 1611) := (wbPartMux(1075) xor i_prn(537)) & (not wbPartMux(1074) xor i_prn(537)) & '1';
    wbMult(1616 downto 1614) := (wbPartMux(1077) xor i_prn(538)) & (not wbPartMux(1076) xor i_prn(538)) & '1';
    wbMult(1619 downto 1617) := (wbPartMux(1079) xor i_prn(539)) & (not wbPartMux(1078) xor i_prn(539)) & '1';
    wbMult(1622 downto 1620) := (wbPartMux(1081) xor i_prn(540)) & (not wbPartMux(1080) xor i_prn(540)) & '1';
    wbMult(1625 downto 1623) := (wbPartMux(1083) xor i_prn(541)) & (not wbPartMux(1082) xor i_prn(541)) & '1';
    wbMult(1628 downto 1626) := (wbPartMux(1085) xor i_prn(542)) & (not wbPartMux(1084) xor i_prn(542)) & '1';
    wbMult(1631 downto 1629) := (wbPartMux(1087) xor i_prn(543)) & (not wbPartMux(1086) xor i_prn(543)) & '1';
    wbMult(1634 downto 1632) := (wbPartMux(1089) xor i_prn(544)) & (not wbPartMux(1088) xor i_prn(544)) & '1';
    wbMult(1637 downto 1635) := (wbPartMux(1091) xor i_prn(545)) & (not wbPartMux(1090) xor i_prn(545)) & '1';
    wbMult(1640 downto 1638) := (wbPartMux(1093) xor i_prn(546)) & (not wbPartMux(1092) xor i_prn(546)) & '1';
    wbMult(1643 downto 1641) := (wbPartMux(1095) xor i_prn(547)) & (not wbPartMux(1094) xor i_prn(547)) & '1';
    wbMult(1646 downto 1644) := (wbPartMux(1097) xor i_prn(548)) & (not wbPartMux(1096) xor i_prn(548)) & '1';
    wbMult(1649 downto 1647) := (wbPartMux(1099) xor i_prn(549)) & (not wbPartMux(1098) xor i_prn(549)) & '1';
    wbMult(1652 downto 1650) := (wbPartMux(1101) xor i_prn(550)) & (not wbPartMux(1100) xor i_prn(550)) & '1';
    wbMult(1655 downto 1653) := (wbPartMux(1103) xor i_prn(551)) & (not wbPartMux(1102) xor i_prn(551)) & '1';
    wbMult(1658 downto 1656) := (wbPartMux(1105) xor i_prn(552)) & (not wbPartMux(1104) xor i_prn(552)) & '1';
    wbMult(1661 downto 1659) := (wbPartMux(1107) xor i_prn(553)) & (not wbPartMux(1106) xor i_prn(553)) & '1';
    wbMult(1664 downto 1662) := (wbPartMux(1109) xor i_prn(554)) & (not wbPartMux(1108) xor i_prn(554)) & '1';
    wbMult(1667 downto 1665) := (wbPartMux(1111) xor i_prn(555)) & (not wbPartMux(1110) xor i_prn(555)) & '1';
    wbMult(1670 downto 1668) := (wbPartMux(1113) xor i_prn(556)) & (not wbPartMux(1112) xor i_prn(556)) & '1';
    wbMult(1673 downto 1671) := (wbPartMux(1115) xor i_prn(557)) & (not wbPartMux(1114) xor i_prn(557)) & '1';
    wbMult(1676 downto 1674) := (wbPartMux(1117) xor i_prn(558)) & (not wbPartMux(1116) xor i_prn(558)) & '1';
    wbMult(1679 downto 1677) := (wbPartMux(1119) xor i_prn(559)) & (not wbPartMux(1118) xor i_prn(559)) & '1';
    wbMult(1682 downto 1680) := (wbPartMux(1121) xor i_prn(560)) & (not wbPartMux(1120) xor i_prn(560)) & '1';
    wbMult(1685 downto 1683) := (wbPartMux(1123) xor i_prn(561)) & (not wbPartMux(1122) xor i_prn(561)) & '1';
    wbMult(1688 downto 1686) := (wbPartMux(1125) xor i_prn(562)) & (not wbPartMux(1124) xor i_prn(562)) & '1';
    wbMult(1691 downto 1689) := (wbPartMux(1127) xor i_prn(563)) & (not wbPartMux(1126) xor i_prn(563)) & '1';
    wbMult(1694 downto 1692) := (wbPartMux(1129) xor i_prn(564)) & (not wbPartMux(1128) xor i_prn(564)) & '1';
    wbMult(1697 downto 1695) := (wbPartMux(1131) xor i_prn(565)) & (not wbPartMux(1130) xor i_prn(565)) & '1';
    wbMult(1700 downto 1698) := (wbPartMux(1133) xor i_prn(566)) & (not wbPartMux(1132) xor i_prn(566)) & '1';
    wbMult(1703 downto 1701) := (wbPartMux(1135) xor i_prn(567)) & (not wbPartMux(1134) xor i_prn(567)) & '1';
    wbMult(1706 downto 1704) := (wbPartMux(1137) xor i_prn(568)) & (not wbPartMux(1136) xor i_prn(568)) & '1';
    wbMult(1709 downto 1707) := (wbPartMux(1139) xor i_prn(569)) & (not wbPartMux(1138) xor i_prn(569)) & '1';
    wbMult(1712 downto 1710) := (wbPartMux(1141) xor i_prn(570)) & (not wbPartMux(1140) xor i_prn(570)) & '1';
    wbMult(1715 downto 1713) := (wbPartMux(1143) xor i_prn(571)) & (not wbPartMux(1142) xor i_prn(571)) & '1';
    wbMult(1718 downto 1716) := (wbPartMux(1145) xor i_prn(572)) & (not wbPartMux(1144) xor i_prn(572)) & '1';
    wbMult(1721 downto 1719) := (wbPartMux(1147) xor i_prn(573)) & (not wbPartMux(1146) xor i_prn(573)) & '1';
    wbMult(1724 downto 1722) := (wbPartMux(1149) xor i_prn(574)) & (not wbPartMux(1148) xor i_prn(574)) & '1';
    wbMult(1727 downto 1725) := (wbPartMux(1151) xor i_prn(575)) & (not wbPartMux(1150) xor i_prn(575)) & '1';
    wbMult(1730 downto 1728) := (wbPartMux(1153) xor i_prn(576)) & (not wbPartMux(1152) xor i_prn(576)) & '1';
    wbMult(1733 downto 1731) := (wbPartMux(1155) xor i_prn(577)) & (not wbPartMux(1154) xor i_prn(577)) & '1';
    wbMult(1736 downto 1734) := (wbPartMux(1157) xor i_prn(578)) & (not wbPartMux(1156) xor i_prn(578)) & '1';
    wbMult(1739 downto 1737) := (wbPartMux(1159) xor i_prn(579)) & (not wbPartMux(1158) xor i_prn(579)) & '1';
    wbMult(1742 downto 1740) := (wbPartMux(1161) xor i_prn(580)) & (not wbPartMux(1160) xor i_prn(580)) & '1';
    wbMult(1745 downto 1743) := (wbPartMux(1163) xor i_prn(581)) & (not wbPartMux(1162) xor i_prn(581)) & '1';
    wbMult(1748 downto 1746) := (wbPartMux(1165) xor i_prn(582)) & (not wbPartMux(1164) xor i_prn(582)) & '1';
    wbMult(1751 downto 1749) := (wbPartMux(1167) xor i_prn(583)) & (not wbPartMux(1166) xor i_prn(583)) & '1';
    wbMult(1754 downto 1752) := (wbPartMux(1169) xor i_prn(584)) & (not wbPartMux(1168) xor i_prn(584)) & '1';
    wbMult(1757 downto 1755) := (wbPartMux(1171) xor i_prn(585)) & (not wbPartMux(1170) xor i_prn(585)) & '1';
    wbMult(1760 downto 1758) := (wbPartMux(1173) xor i_prn(586)) & (not wbPartMux(1172) xor i_prn(586)) & '1';
    wbMult(1763 downto 1761) := (wbPartMux(1175) xor i_prn(587)) & (not wbPartMux(1174) xor i_prn(587)) & '1';
    wbMult(1766 downto 1764) := (wbPartMux(1177) xor i_prn(588)) & (not wbPartMux(1176) xor i_prn(588)) & '1';
    wbMult(1769 downto 1767) := (wbPartMux(1179) xor i_prn(589)) & (not wbPartMux(1178) xor i_prn(589)) & '1';
    wbMult(1772 downto 1770) := (wbPartMux(1181) xor i_prn(590)) & (not wbPartMux(1180) xor i_prn(590)) & '1';
    wbMult(1775 downto 1773) := (wbPartMux(1183) xor i_prn(591)) & (not wbPartMux(1182) xor i_prn(591)) & '1';
    wbMult(1778 downto 1776) := (wbPartMux(1185) xor i_prn(592)) & (not wbPartMux(1184) xor i_prn(592)) & '1';
    wbMult(1781 downto 1779) := (wbPartMux(1187) xor i_prn(593)) & (not wbPartMux(1186) xor i_prn(593)) & '1';
    wbMult(1784 downto 1782) := (wbPartMux(1189) xor i_prn(594)) & (not wbPartMux(1188) xor i_prn(594)) & '1';
    wbMult(1787 downto 1785) := (wbPartMux(1191) xor i_prn(595)) & (not wbPartMux(1190) xor i_prn(595)) & '1';
    wbMult(1790 downto 1788) := (wbPartMux(1193) xor i_prn(596)) & (not wbPartMux(1192) xor i_prn(596)) & '1';
    wbMult(1793 downto 1791) := (wbPartMux(1195) xor i_prn(597)) & (not wbPartMux(1194) xor i_prn(597)) & '1';
    wbMult(1796 downto 1794) := (wbPartMux(1197) xor i_prn(598)) & (not wbPartMux(1196) xor i_prn(598)) & '1';
    wbMult(1799 downto 1797) := (wbPartMux(1199) xor i_prn(599)) & (not wbPartMux(1198) xor i_prn(599)) & '1';
    wbMult(1802 downto 1800) := (wbPartMux(1201) xor i_prn(600)) & (not wbPartMux(1200) xor i_prn(600)) & '1';
    wbMult(1805 downto 1803) := (wbPartMux(1203) xor i_prn(601)) & (not wbPartMux(1202) xor i_prn(601)) & '1';
    wbMult(1808 downto 1806) := (wbPartMux(1205) xor i_prn(602)) & (not wbPartMux(1204) xor i_prn(602)) & '1';
    wbMult(1811 downto 1809) := (wbPartMux(1207) xor i_prn(603)) & (not wbPartMux(1206) xor i_prn(603)) & '1';
    wbMult(1814 downto 1812) := (wbPartMux(1209) xor i_prn(604)) & (not wbPartMux(1208) xor i_prn(604)) & '1';
    wbMult(1817 downto 1815) := (wbPartMux(1211) xor i_prn(605)) & (not wbPartMux(1210) xor i_prn(605)) & '1';
    wbMult(1820 downto 1818) := (wbPartMux(1213) xor i_prn(606)) & (not wbPartMux(1212) xor i_prn(606)) & '1';
    wbMult(1823 downto 1821) := (wbPartMux(1215) xor i_prn(607)) & (not wbPartMux(1214) xor i_prn(607)) & '1';
    wbMult(1826 downto 1824) := (wbPartMux(1217) xor i_prn(608)) & (not wbPartMux(1216) xor i_prn(608)) & '1';
    wbMult(1829 downto 1827) := (wbPartMux(1219) xor i_prn(609)) & (not wbPartMux(1218) xor i_prn(609)) & '1';
    wbMult(1832 downto 1830) := (wbPartMux(1221) xor i_prn(610)) & (not wbPartMux(1220) xor i_prn(610)) & '1';
    wbMult(1835 downto 1833) := (wbPartMux(1223) xor i_prn(611)) & (not wbPartMux(1222) xor i_prn(611)) & '1';
    wbMult(1838 downto 1836) := (wbPartMux(1225) xor i_prn(612)) & (not wbPartMux(1224) xor i_prn(612)) & '1';
    wbMult(1841 downto 1839) := (wbPartMux(1227) xor i_prn(613)) & (not wbPartMux(1226) xor i_prn(613)) & '1';
    wbMult(1844 downto 1842) := (wbPartMux(1229) xor i_prn(614)) & (not wbPartMux(1228) xor i_prn(614)) & '1';
    wbMult(1847 downto 1845) := (wbPartMux(1231) xor i_prn(615)) & (not wbPartMux(1230) xor i_prn(615)) & '1';
    wbMult(1850 downto 1848) := (wbPartMux(1233) xor i_prn(616)) & (not wbPartMux(1232) xor i_prn(616)) & '1';
    wbMult(1853 downto 1851) := (wbPartMux(1235) xor i_prn(617)) & (not wbPartMux(1234) xor i_prn(617)) & '1';
    wbMult(1856 downto 1854) := (wbPartMux(1237) xor i_prn(618)) & (not wbPartMux(1236) xor i_prn(618)) & '1';
    wbMult(1859 downto 1857) := (wbPartMux(1239) xor i_prn(619)) & (not wbPartMux(1238) xor i_prn(619)) & '1';
    wbMult(1862 downto 1860) := (wbPartMux(1241) xor i_prn(620)) & (not wbPartMux(1240) xor i_prn(620)) & '1';
    wbMult(1865 downto 1863) := (wbPartMux(1243) xor i_prn(621)) & (not wbPartMux(1242) xor i_prn(621)) & '1';
    wbMult(1868 downto 1866) := (wbPartMux(1245) xor i_prn(622)) & (not wbPartMux(1244) xor i_prn(622)) & '1';
    wbMult(1871 downto 1869) := (wbPartMux(1247) xor i_prn(623)) & (not wbPartMux(1246) xor i_prn(623)) & '1';
    wbMult(1874 downto 1872) := (wbPartMux(1249) xor i_prn(624)) & (not wbPartMux(1248) xor i_prn(624)) & '1';
    wbMult(1877 downto 1875) := (wbPartMux(1251) xor i_prn(625)) & (not wbPartMux(1250) xor i_prn(625)) & '1';
    wbMult(1880 downto 1878) := (wbPartMux(1253) xor i_prn(626)) & (not wbPartMux(1252) xor i_prn(626)) & '1';
    wbMult(1883 downto 1881) := (wbPartMux(1255) xor i_prn(627)) & (not wbPartMux(1254) xor i_prn(627)) & '1';
    wbMult(1886 downto 1884) := (wbPartMux(1257) xor i_prn(628)) & (not wbPartMux(1256) xor i_prn(628)) & '1';
    wbMult(1889 downto 1887) := (wbPartMux(1259) xor i_prn(629)) & (not wbPartMux(1258) xor i_prn(629)) & '1';
    wbMult(1892 downto 1890) := (wbPartMux(1261) xor i_prn(630)) & (not wbPartMux(1260) xor i_prn(630)) & '1';
    wbMult(1895 downto 1893) := (wbPartMux(1263) xor i_prn(631)) & (not wbPartMux(1262) xor i_prn(631)) & '1';
    wbMult(1898 downto 1896) := (wbPartMux(1265) xor i_prn(632)) & (not wbPartMux(1264) xor i_prn(632)) & '1';
    wbMult(1901 downto 1899) := (wbPartMux(1267) xor i_prn(633)) & (not wbPartMux(1266) xor i_prn(633)) & '1';
    wbMult(1904 downto 1902) := (wbPartMux(1269) xor i_prn(634)) & (not wbPartMux(1268) xor i_prn(634)) & '1';
    wbMult(1907 downto 1905) := (wbPartMux(1271) xor i_prn(635)) & (not wbPartMux(1270) xor i_prn(635)) & '1';
    wbMult(1910 downto 1908) := (wbPartMux(1273) xor i_prn(636)) & (not wbPartMux(1272) xor i_prn(636)) & '1';
    wbMult(1913 downto 1911) := (wbPartMux(1275) xor i_prn(637)) & (not wbPartMux(1274) xor i_prn(637)) & '1';
    wbMult(1916 downto 1914) := (wbPartMux(1277) xor i_prn(638)) & (not wbPartMux(1276) xor i_prn(638)) & '1';
    wbMult(1919 downto 1917) := (wbPartMux(1279) xor i_prn(639)) & (not wbPartMux(1278) xor i_prn(639)) & '1';
    wbMult(1922 downto 1920) := (wbPartMux(1281) xor i_prn(640)) & (not wbPartMux(1280) xor i_prn(640)) & '1';
    wbMult(1925 downto 1923) := (wbPartMux(1283) xor i_prn(641)) & (not wbPartMux(1282) xor i_prn(641)) & '1';
    wbMult(1928 downto 1926) := (wbPartMux(1285) xor i_prn(642)) & (not wbPartMux(1284) xor i_prn(642)) & '1';
    wbMult(1931 downto 1929) := (wbPartMux(1287) xor i_prn(643)) & (not wbPartMux(1286) xor i_prn(643)) & '1';
    wbMult(1934 downto 1932) := (wbPartMux(1289) xor i_prn(644)) & (not wbPartMux(1288) xor i_prn(644)) & '1';
    wbMult(1937 downto 1935) := (wbPartMux(1291) xor i_prn(645)) & (not wbPartMux(1290) xor i_prn(645)) & '1';
    wbMult(1940 downto 1938) := (wbPartMux(1293) xor i_prn(646)) & (not wbPartMux(1292) xor i_prn(646)) & '1';
    wbMult(1943 downto 1941) := (wbPartMux(1295) xor i_prn(647)) & (not wbPartMux(1294) xor i_prn(647)) & '1';
    wbMult(1946 downto 1944) := (wbPartMux(1297) xor i_prn(648)) & (not wbPartMux(1296) xor i_prn(648)) & '1';
    wbMult(1949 downto 1947) := (wbPartMux(1299) xor i_prn(649)) & (not wbPartMux(1298) xor i_prn(649)) & '1';
    wbMult(1952 downto 1950) := (wbPartMux(1301) xor i_prn(650)) & (not wbPartMux(1300) xor i_prn(650)) & '1';
    wbMult(1955 downto 1953) := (wbPartMux(1303) xor i_prn(651)) & (not wbPartMux(1302) xor i_prn(651)) & '1';
    wbMult(1958 downto 1956) := (wbPartMux(1305) xor i_prn(652)) & (not wbPartMux(1304) xor i_prn(652)) & '1';
    wbMult(1961 downto 1959) := (wbPartMux(1307) xor i_prn(653)) & (not wbPartMux(1306) xor i_prn(653)) & '1';
    wbMult(1964 downto 1962) := (wbPartMux(1309) xor i_prn(654)) & (not wbPartMux(1308) xor i_prn(654)) & '1';
    wbMult(1967 downto 1965) := (wbPartMux(1311) xor i_prn(655)) & (not wbPartMux(1310) xor i_prn(655)) & '1';
    wbMult(1970 downto 1968) := (wbPartMux(1313) xor i_prn(656)) & (not wbPartMux(1312) xor i_prn(656)) & '1';
    wbMult(1973 downto 1971) := (wbPartMux(1315) xor i_prn(657)) & (not wbPartMux(1314) xor i_prn(657)) & '1';
    wbMult(1976 downto 1974) := (wbPartMux(1317) xor i_prn(658)) & (not wbPartMux(1316) xor i_prn(658)) & '1';
    wbMult(1979 downto 1977) := (wbPartMux(1319) xor i_prn(659)) & (not wbPartMux(1318) xor i_prn(659)) & '1';
    wbMult(1982 downto 1980) := (wbPartMux(1321) xor i_prn(660)) & (not wbPartMux(1320) xor i_prn(660)) & '1';
    wbMult(1985 downto 1983) := (wbPartMux(1323) xor i_prn(661)) & (not wbPartMux(1322) xor i_prn(661)) & '1';
    wbMult(1988 downto 1986) := (wbPartMux(1325) xor i_prn(662)) & (not wbPartMux(1324) xor i_prn(662)) & '1';
    wbMult(1991 downto 1989) := (wbPartMux(1327) xor i_prn(663)) & (not wbPartMux(1326) xor i_prn(663)) & '1';
    wbMult(1994 downto 1992) := (wbPartMux(1329) xor i_prn(664)) & (not wbPartMux(1328) xor i_prn(664)) & '1';
    wbMult(1997 downto 1995) := (wbPartMux(1331) xor i_prn(665)) & (not wbPartMux(1330) xor i_prn(665)) & '1';
    wbMult(2000 downto 1998) := (wbPartMux(1333) xor i_prn(666)) & (not wbPartMux(1332) xor i_prn(666)) & '1';
    wbMult(2003 downto 2001) := (wbPartMux(1335) xor i_prn(667)) & (not wbPartMux(1334) xor i_prn(667)) & '1';
    wbMult(2006 downto 2004) := (wbPartMux(1337) xor i_prn(668)) & (not wbPartMux(1336) xor i_prn(668)) & '1';
    wbMult(2009 downto 2007) := (wbPartMux(1339) xor i_prn(669)) & (not wbPartMux(1338) xor i_prn(669)) & '1';
    wbMult(2012 downto 2010) := (wbPartMux(1341) xor i_prn(670)) & (not wbPartMux(1340) xor i_prn(670)) & '1';
    wbMult(2015 downto 2013) := (wbPartMux(1343) xor i_prn(671)) & (not wbPartMux(1342) xor i_prn(671)) & '1';
    wbMult(2018 downto 2016) := (wbPartMux(1345) xor i_prn(672)) & (not wbPartMux(1344) xor i_prn(672)) & '1';
    wbMult(2021 downto 2019) := (wbPartMux(1347) xor i_prn(673)) & (not wbPartMux(1346) xor i_prn(673)) & '1';
    wbMult(2024 downto 2022) := (wbPartMux(1349) xor i_prn(674)) & (not wbPartMux(1348) xor i_prn(674)) & '1';
    wbMult(2027 downto 2025) := (wbPartMux(1351) xor i_prn(675)) & (not wbPartMux(1350) xor i_prn(675)) & '1';
    wbMult(2030 downto 2028) := (wbPartMux(1353) xor i_prn(676)) & (not wbPartMux(1352) xor i_prn(676)) & '1';
    wbMult(2033 downto 2031) := (wbPartMux(1355) xor i_prn(677)) & (not wbPartMux(1354) xor i_prn(677)) & '1';
    wbMult(2036 downto 2034) := (wbPartMux(1357) xor i_prn(678)) & (not wbPartMux(1356) xor i_prn(678)) & '1';
    wbMult(2039 downto 2037) := (wbPartMux(1359) xor i_prn(679)) & (not wbPartMux(1358) xor i_prn(679)) & '1';
    wbMult(2042 downto 2040) := (wbPartMux(1361) xor i_prn(680)) & (not wbPartMux(1360) xor i_prn(680)) & '1';
    wbMult(2045 downto 2043) := (wbPartMux(1363) xor i_prn(681)) & (not wbPartMux(1362) xor i_prn(681)) & '1';
    wbMult(2048 downto 2046) := (wbPartMux(1365) xor i_prn(682)) & (not wbPartMux(1364) xor i_prn(682)) & '1';
    wbMult(2051 downto 2049) := (wbPartMux(1367) xor i_prn(683)) & (not wbPartMux(1366) xor i_prn(683)) & '1';
    wbMult(2054 downto 2052) := (wbPartMux(1369) xor i_prn(684)) & (not wbPartMux(1368) xor i_prn(684)) & '1';
    wbMult(2057 downto 2055) := (wbPartMux(1371) xor i_prn(685)) & (not wbPartMux(1370) xor i_prn(685)) & '1';
    wbMult(2060 downto 2058) := (wbPartMux(1373) xor i_prn(686)) & (not wbPartMux(1372) xor i_prn(686)) & '1';
    wbMult(2063 downto 2061) := (wbPartMux(1375) xor i_prn(687)) & (not wbPartMux(1374) xor i_prn(687)) & '1';
    wbMult(2066 downto 2064) := (wbPartMux(1377) xor i_prn(688)) & (not wbPartMux(1376) xor i_prn(688)) & '1';
    wbMult(2069 downto 2067) := (wbPartMux(1379) xor i_prn(689)) & (not wbPartMux(1378) xor i_prn(689)) & '1';
    wbMult(2072 downto 2070) := (wbPartMux(1381) xor i_prn(690)) & (not wbPartMux(1380) xor i_prn(690)) & '1';
    wbMult(2075 downto 2073) := (wbPartMux(1383) xor i_prn(691)) & (not wbPartMux(1382) xor i_prn(691)) & '1';
    wbMult(2078 downto 2076) := (wbPartMux(1385) xor i_prn(692)) & (not wbPartMux(1384) xor i_prn(692)) & '1';
    wbMult(2081 downto 2079) := (wbPartMux(1387) xor i_prn(693)) & (not wbPartMux(1386) xor i_prn(693)) & '1';
    wbMult(2084 downto 2082) := (wbPartMux(1389) xor i_prn(694)) & (not wbPartMux(1388) xor i_prn(694)) & '1';
    wbMult(2087 downto 2085) := (wbPartMux(1391) xor i_prn(695)) & (not wbPartMux(1390) xor i_prn(695)) & '1';
    wbMult(2090 downto 2088) := (wbPartMux(1393) xor i_prn(696)) & (not wbPartMux(1392) xor i_prn(696)) & '1';
    wbMult(2093 downto 2091) := (wbPartMux(1395) xor i_prn(697)) & (not wbPartMux(1394) xor i_prn(697)) & '1';
    wbMult(2096 downto 2094) := (wbPartMux(1397) xor i_prn(698)) & (not wbPartMux(1396) xor i_prn(698)) & '1';
    wbMult(2099 downto 2097) := (wbPartMux(1399) xor i_prn(699)) & (not wbPartMux(1398) xor i_prn(699)) & '1';
    wbMult(2102 downto 2100) := (wbPartMux(1401) xor i_prn(700)) & (not wbPartMux(1400) xor i_prn(700)) & '1';
    wbMult(2105 downto 2103) := (wbPartMux(1403) xor i_prn(701)) & (not wbPartMux(1402) xor i_prn(701)) & '1';
    wbMult(2108 downto 2106) := (wbPartMux(1405) xor i_prn(702)) & (not wbPartMux(1404) xor i_prn(702)) & '1';
    wbMult(2111 downto 2109) := (wbPartMux(1407) xor i_prn(703)) & (not wbPartMux(1406) xor i_prn(703)) & '1';
    wbMult(2114 downto 2112) := (wbPartMux(1409) xor i_prn(704)) & (not wbPartMux(1408) xor i_prn(704)) & '1';
    wbMult(2117 downto 2115) := (wbPartMux(1411) xor i_prn(705)) & (not wbPartMux(1410) xor i_prn(705)) & '1';
    wbMult(2120 downto 2118) := (wbPartMux(1413) xor i_prn(706)) & (not wbPartMux(1412) xor i_prn(706)) & '1';
    wbMult(2123 downto 2121) := (wbPartMux(1415) xor i_prn(707)) & (not wbPartMux(1414) xor i_prn(707)) & '1';
    wbMult(2126 downto 2124) := (wbPartMux(1417) xor i_prn(708)) & (not wbPartMux(1416) xor i_prn(708)) & '1';
    wbMult(2129 downto 2127) := (wbPartMux(1419) xor i_prn(709)) & (not wbPartMux(1418) xor i_prn(709)) & '1';
    wbMult(2132 downto 2130) := (wbPartMux(1421) xor i_prn(710)) & (not wbPartMux(1420) xor i_prn(710)) & '1';
    wbMult(2135 downto 2133) := (wbPartMux(1423) xor i_prn(711)) & (not wbPartMux(1422) xor i_prn(711)) & '1';
    wbMult(2138 downto 2136) := (wbPartMux(1425) xor i_prn(712)) & (not wbPartMux(1424) xor i_prn(712)) & '1';
    wbMult(2141 downto 2139) := (wbPartMux(1427) xor i_prn(713)) & (not wbPartMux(1426) xor i_prn(713)) & '1';
    wbMult(2144 downto 2142) := (wbPartMux(1429) xor i_prn(714)) & (not wbPartMux(1428) xor i_prn(714)) & '1';
    wbMult(2147 downto 2145) := (wbPartMux(1431) xor i_prn(715)) & (not wbPartMux(1430) xor i_prn(715)) & '1';
    wbMult(2150 downto 2148) := (wbPartMux(1433) xor i_prn(716)) & (not wbPartMux(1432) xor i_prn(716)) & '1';
    wbMult(2153 downto 2151) := (wbPartMux(1435) xor i_prn(717)) & (not wbPartMux(1434) xor i_prn(717)) & '1';
    wbMult(2156 downto 2154) := (wbPartMux(1437) xor i_prn(718)) & (not wbPartMux(1436) xor i_prn(718)) & '1';
    wbMult(2159 downto 2157) := (wbPartMux(1439) xor i_prn(719)) & (not wbPartMux(1438) xor i_prn(719)) & '1';
    wbMult(2162 downto 2160) := (wbPartMux(1441) xor i_prn(720)) & (not wbPartMux(1440) xor i_prn(720)) & '1';
    wbMult(2165 downto 2163) := (wbPartMux(1443) xor i_prn(721)) & (not wbPartMux(1442) xor i_prn(721)) & '1';
    wbMult(2168 downto 2166) := (wbPartMux(1445) xor i_prn(722)) & (not wbPartMux(1444) xor i_prn(722)) & '1';
    wbMult(2171 downto 2169) := (wbPartMux(1447) xor i_prn(723)) & (not wbPartMux(1446) xor i_prn(723)) & '1';
    wbMult(2174 downto 2172) := (wbPartMux(1449) xor i_prn(724)) & (not wbPartMux(1448) xor i_prn(724)) & '1';
    wbMult(2177 downto 2175) := (wbPartMux(1451) xor i_prn(725)) & (not wbPartMux(1450) xor i_prn(725)) & '1';
    wbMult(2180 downto 2178) := (wbPartMux(1453) xor i_prn(726)) & (not wbPartMux(1452) xor i_prn(726)) & '1';
    wbMult(2183 downto 2181) := (wbPartMux(1455) xor i_prn(727)) & (not wbPartMux(1454) xor i_prn(727)) & '1';
    wbMult(2186 downto 2184) := (wbPartMux(1457) xor i_prn(728)) & (not wbPartMux(1456) xor i_prn(728)) & '1';
    wbMult(2189 downto 2187) := (wbPartMux(1459) xor i_prn(729)) & (not wbPartMux(1458) xor i_prn(729)) & '1';
    wbMult(2192 downto 2190) := (wbPartMux(1461) xor i_prn(730)) & (not wbPartMux(1460) xor i_prn(730)) & '1';
    wbMult(2195 downto 2193) := (wbPartMux(1463) xor i_prn(731)) & (not wbPartMux(1462) xor i_prn(731)) & '1';
    wbMult(2198 downto 2196) := (wbPartMux(1465) xor i_prn(732)) & (not wbPartMux(1464) xor i_prn(732)) & '1';
    wbMult(2201 downto 2199) := (wbPartMux(1467) xor i_prn(733)) & (not wbPartMux(1466) xor i_prn(733)) & '1';
    wbMult(2204 downto 2202) := (wbPartMux(1469) xor i_prn(734)) & (not wbPartMux(1468) xor i_prn(734)) & '1';
    wbMult(2207 downto 2205) := (wbPartMux(1471) xor i_prn(735)) & (not wbPartMux(1470) xor i_prn(735)) & '1';
    wbMult(2210 downto 2208) := (wbPartMux(1473) xor i_prn(736)) & (not wbPartMux(1472) xor i_prn(736)) & '1';
    wbMult(2213 downto 2211) := (wbPartMux(1475) xor i_prn(737)) & (not wbPartMux(1474) xor i_prn(737)) & '1';
    wbMult(2216 downto 2214) := (wbPartMux(1477) xor i_prn(738)) & (not wbPartMux(1476) xor i_prn(738)) & '1';
    wbMult(2219 downto 2217) := (wbPartMux(1479) xor i_prn(739)) & (not wbPartMux(1478) xor i_prn(739)) & '1';
    wbMult(2222 downto 2220) := (wbPartMux(1481) xor i_prn(740)) & (not wbPartMux(1480) xor i_prn(740)) & '1';
    wbMult(2225 downto 2223) := (wbPartMux(1483) xor i_prn(741)) & (not wbPartMux(1482) xor i_prn(741)) & '1';
    wbMult(2228 downto 2226) := (wbPartMux(1485) xor i_prn(742)) & (not wbPartMux(1484) xor i_prn(742)) & '1';
    wbMult(2231 downto 2229) := (wbPartMux(1487) xor i_prn(743)) & (not wbPartMux(1486) xor i_prn(743)) & '1';
    wbMult(2234 downto 2232) := (wbPartMux(1489) xor i_prn(744)) & (not wbPartMux(1488) xor i_prn(744)) & '1';
    wbMult(2237 downto 2235) := (wbPartMux(1491) xor i_prn(745)) & (not wbPartMux(1490) xor i_prn(745)) & '1';
    wbMult(2240 downto 2238) := (wbPartMux(1493) xor i_prn(746)) & (not wbPartMux(1492) xor i_prn(746)) & '1';
    wbMult(2243 downto 2241) := (wbPartMux(1495) xor i_prn(747)) & (not wbPartMux(1494) xor i_prn(747)) & '1';
    wbMult(2246 downto 2244) := (wbPartMux(1497) xor i_prn(748)) & (not wbPartMux(1496) xor i_prn(748)) & '1';
    wbMult(2249 downto 2247) := (wbPartMux(1499) xor i_prn(749)) & (not wbPartMux(1498) xor i_prn(749)) & '1';
    wbMult(2252 downto 2250) := (wbPartMux(1501) xor i_prn(750)) & (not wbPartMux(1500) xor i_prn(750)) & '1';
    wbMult(2255 downto 2253) := (wbPartMux(1503) xor i_prn(751)) & (not wbPartMux(1502) xor i_prn(751)) & '1';
    wbMult(2258 downto 2256) := (wbPartMux(1505) xor i_prn(752)) & (not wbPartMux(1504) xor i_prn(752)) & '1';
    wbMult(2261 downto 2259) := (wbPartMux(1507) xor i_prn(753)) & (not wbPartMux(1506) xor i_prn(753)) & '1';
    wbMult(2264 downto 2262) := (wbPartMux(1509) xor i_prn(754)) & (not wbPartMux(1508) xor i_prn(754)) & '1';
    wbMult(2267 downto 2265) := (wbPartMux(1511) xor i_prn(755)) & (not wbPartMux(1510) xor i_prn(755)) & '1';
    wbMult(2270 downto 2268) := (wbPartMux(1513) xor i_prn(756)) & (not wbPartMux(1512) xor i_prn(756)) & '1';
    wbMult(2273 downto 2271) := (wbPartMux(1515) xor i_prn(757)) & (not wbPartMux(1514) xor i_prn(757)) & '1';
    wbMult(2276 downto 2274) := (wbPartMux(1517) xor i_prn(758)) & (not wbPartMux(1516) xor i_prn(758)) & '1';
    wbMult(2279 downto 2277) := (wbPartMux(1519) xor i_prn(759)) & (not wbPartMux(1518) xor i_prn(759)) & '1';
    wbMult(2282 downto 2280) := (wbPartMux(1521) xor i_prn(760)) & (not wbPartMux(1520) xor i_prn(760)) & '1';
    wbMult(2285 downto 2283) := (wbPartMux(1523) xor i_prn(761)) & (not wbPartMux(1522) xor i_prn(761)) & '1';
    wbMult(2288 downto 2286) := (wbPartMux(1525) xor i_prn(762)) & (not wbPartMux(1524) xor i_prn(762)) & '1';
    wbMult(2291 downto 2289) := (wbPartMux(1527) xor i_prn(763)) & (not wbPartMux(1526) xor i_prn(763)) & '1';
    wbMult(2294 downto 2292) := (wbPartMux(1529) xor i_prn(764)) & (not wbPartMux(1528) xor i_prn(764)) & '1';
    wbMult(2297 downto 2295) := (wbPartMux(1531) xor i_prn(765)) & (not wbPartMux(1530) xor i_prn(765)) & '1';
    wbMult(2300 downto 2298) := (wbPartMux(1533) xor i_prn(766)) & (not wbPartMux(1532) xor i_prn(766)) & '1';
    wbMult(2303 downto 2301) := (wbPartMux(1535) xor i_prn(767)) & (not wbPartMux(1534) xor i_prn(767)) & '1';
    wbMult(2306 downto 2304) := (wbPartMux(1537) xor i_prn(768)) & (not wbPartMux(1536) xor i_prn(768)) & '1';
    wbMult(2309 downto 2307) := (wbPartMux(1539) xor i_prn(769)) & (not wbPartMux(1538) xor i_prn(769)) & '1';
    wbMult(2312 downto 2310) := (wbPartMux(1541) xor i_prn(770)) & (not wbPartMux(1540) xor i_prn(770)) & '1';
    wbMult(2315 downto 2313) := (wbPartMux(1543) xor i_prn(771)) & (not wbPartMux(1542) xor i_prn(771)) & '1';
    wbMult(2318 downto 2316) := (wbPartMux(1545) xor i_prn(772)) & (not wbPartMux(1544) xor i_prn(772)) & '1';
    wbMult(2321 downto 2319) := (wbPartMux(1547) xor i_prn(773)) & (not wbPartMux(1546) xor i_prn(773)) & '1';
    wbMult(2324 downto 2322) := (wbPartMux(1549) xor i_prn(774)) & (not wbPartMux(1548) xor i_prn(774)) & '1';
    wbMult(2327 downto 2325) := (wbPartMux(1551) xor i_prn(775)) & (not wbPartMux(1550) xor i_prn(775)) & '1';
    wbMult(2330 downto 2328) := (wbPartMux(1553) xor i_prn(776)) & (not wbPartMux(1552) xor i_prn(776)) & '1';
    wbMult(2333 downto 2331) := (wbPartMux(1555) xor i_prn(777)) & (not wbPartMux(1554) xor i_prn(777)) & '1';
    wbMult(2336 downto 2334) := (wbPartMux(1557) xor i_prn(778)) & (not wbPartMux(1556) xor i_prn(778)) & '1';
    wbMult(2339 downto 2337) := (wbPartMux(1559) xor i_prn(779)) & (not wbPartMux(1558) xor i_prn(779)) & '1';
    wbMult(2342 downto 2340) := (wbPartMux(1561) xor i_prn(780)) & (not wbPartMux(1560) xor i_prn(780)) & '1';
    wbMult(2345 downto 2343) := (wbPartMux(1563) xor i_prn(781)) & (not wbPartMux(1562) xor i_prn(781)) & '1';
    wbMult(2348 downto 2346) := (wbPartMux(1565) xor i_prn(782)) & (not wbPartMux(1564) xor i_prn(782)) & '1';
    wbMult(2351 downto 2349) := (wbPartMux(1567) xor i_prn(783)) & (not wbPartMux(1566) xor i_prn(783)) & '1';
    wbMult(2354 downto 2352) := (wbPartMux(1569) xor i_prn(784)) & (not wbPartMux(1568) xor i_prn(784)) & '1';
    wbMult(2357 downto 2355) := (wbPartMux(1571) xor i_prn(785)) & (not wbPartMux(1570) xor i_prn(785)) & '1';
    wbMult(2360 downto 2358) := (wbPartMux(1573) xor i_prn(786)) & (not wbPartMux(1572) xor i_prn(786)) & '1';
    wbMult(2363 downto 2361) := (wbPartMux(1575) xor i_prn(787)) & (not wbPartMux(1574) xor i_prn(787)) & '1';
    wbMult(2366 downto 2364) := (wbPartMux(1577) xor i_prn(788)) & (not wbPartMux(1576) xor i_prn(788)) & '1';
    wbMult(2369 downto 2367) := (wbPartMux(1579) xor i_prn(789)) & (not wbPartMux(1578) xor i_prn(789)) & '1';
    wbMult(2372 downto 2370) := (wbPartMux(1581) xor i_prn(790)) & (not wbPartMux(1580) xor i_prn(790)) & '1';
    wbMult(2375 downto 2373) := (wbPartMux(1583) xor i_prn(791)) & (not wbPartMux(1582) xor i_prn(791)) & '1';
    wbMult(2378 downto 2376) := (wbPartMux(1585) xor i_prn(792)) & (not wbPartMux(1584) xor i_prn(792)) & '1';
    wbMult(2381 downto 2379) := (wbPartMux(1587) xor i_prn(793)) & (not wbPartMux(1586) xor i_prn(793)) & '1';
    wbMult(2384 downto 2382) := (wbPartMux(1589) xor i_prn(794)) & (not wbPartMux(1588) xor i_prn(794)) & '1';
    wbMult(2387 downto 2385) := (wbPartMux(1591) xor i_prn(795)) & (not wbPartMux(1590) xor i_prn(795)) & '1';
    wbMult(2390 downto 2388) := (wbPartMux(1593) xor i_prn(796)) & (not wbPartMux(1592) xor i_prn(796)) & '1';
    wbMult(2393 downto 2391) := (wbPartMux(1595) xor i_prn(797)) & (not wbPartMux(1594) xor i_prn(797)) & '1';
    wbMult(2396 downto 2394) := (wbPartMux(1597) xor i_prn(798)) & (not wbPartMux(1596) xor i_prn(798)) & '1';
    wbMult(2399 downto 2397) := (wbPartMux(1599) xor i_prn(799)) & (not wbPartMux(1598) xor i_prn(799)) & '1';
    wbMult(2402 downto 2400) := (wbPartMux(1601) xor i_prn(800)) & (not wbPartMux(1600) xor i_prn(800)) & '1';
    wbMult(2405 downto 2403) := (wbPartMux(1603) xor i_prn(801)) & (not wbPartMux(1602) xor i_prn(801)) & '1';
    wbMult(2408 downto 2406) := (wbPartMux(1605) xor i_prn(802)) & (not wbPartMux(1604) xor i_prn(802)) & '1';
    wbMult(2411 downto 2409) := (wbPartMux(1607) xor i_prn(803)) & (not wbPartMux(1606) xor i_prn(803)) & '1';
    wbMult(2414 downto 2412) := (wbPartMux(1609) xor i_prn(804)) & (not wbPartMux(1608) xor i_prn(804)) & '1';
    wbMult(2417 downto 2415) := (wbPartMux(1611) xor i_prn(805)) & (not wbPartMux(1610) xor i_prn(805)) & '1';
    wbMult(2420 downto 2418) := (wbPartMux(1613) xor i_prn(806)) & (not wbPartMux(1612) xor i_prn(806)) & '1';
    wbMult(2423 downto 2421) := (wbPartMux(1615) xor i_prn(807)) & (not wbPartMux(1614) xor i_prn(807)) & '1';
    wbMult(2426 downto 2424) := (wbPartMux(1617) xor i_prn(808)) & (not wbPartMux(1616) xor i_prn(808)) & '1';
    wbMult(2429 downto 2427) := (wbPartMux(1619) xor i_prn(809)) & (not wbPartMux(1618) xor i_prn(809)) & '1';
    wbMult(2432 downto 2430) := (wbPartMux(1621) xor i_prn(810)) & (not wbPartMux(1620) xor i_prn(810)) & '1';
    wbMult(2435 downto 2433) := (wbPartMux(1623) xor i_prn(811)) & (not wbPartMux(1622) xor i_prn(811)) & '1';
    wbMult(2438 downto 2436) := (wbPartMux(1625) xor i_prn(812)) & (not wbPartMux(1624) xor i_prn(812)) & '1';
    wbMult(2441 downto 2439) := (wbPartMux(1627) xor i_prn(813)) & (not wbPartMux(1626) xor i_prn(813)) & '1';
    wbMult(2444 downto 2442) := (wbPartMux(1629) xor i_prn(814)) & (not wbPartMux(1628) xor i_prn(814)) & '1';
    wbMult(2447 downto 2445) := (wbPartMux(1631) xor i_prn(815)) & (not wbPartMux(1630) xor i_prn(815)) & '1';
    wbMult(2450 downto 2448) := (wbPartMux(1633) xor i_prn(816)) & (not wbPartMux(1632) xor i_prn(816)) & '1';
    wbMult(2453 downto 2451) := (wbPartMux(1635) xor i_prn(817)) & (not wbPartMux(1634) xor i_prn(817)) & '1';
    wbMult(2456 downto 2454) := (wbPartMux(1637) xor i_prn(818)) & (not wbPartMux(1636) xor i_prn(818)) & '1';
    wbMult(2459 downto 2457) := (wbPartMux(1639) xor i_prn(819)) & (not wbPartMux(1638) xor i_prn(819)) & '1';
    wbMult(2462 downto 2460) := (wbPartMux(1641) xor i_prn(820)) & (not wbPartMux(1640) xor i_prn(820)) & '1';
    wbMult(2465 downto 2463) := (wbPartMux(1643) xor i_prn(821)) & (not wbPartMux(1642) xor i_prn(821)) & '1';
    wbMult(2468 downto 2466) := (wbPartMux(1645) xor i_prn(822)) & (not wbPartMux(1644) xor i_prn(822)) & '1';
    wbMult(2471 downto 2469) := (wbPartMux(1647) xor i_prn(823)) & (not wbPartMux(1646) xor i_prn(823)) & '1';
    wbMult(2474 downto 2472) := (wbPartMux(1649) xor i_prn(824)) & (not wbPartMux(1648) xor i_prn(824)) & '1';
    wbMult(2477 downto 2475) := (wbPartMux(1651) xor i_prn(825)) & (not wbPartMux(1650) xor i_prn(825)) & '1';
    wbMult(2480 downto 2478) := (wbPartMux(1653) xor i_prn(826)) & (not wbPartMux(1652) xor i_prn(826)) & '1';
    wbMult(2483 downto 2481) := (wbPartMux(1655) xor i_prn(827)) & (not wbPartMux(1654) xor i_prn(827)) & '1';
    wbMult(2486 downto 2484) := (wbPartMux(1657) xor i_prn(828)) & (not wbPartMux(1656) xor i_prn(828)) & '1';
    wbMult(2489 downto 2487) := (wbPartMux(1659) xor i_prn(829)) & (not wbPartMux(1658) xor i_prn(829)) & '1';
    wbMult(2492 downto 2490) := (wbPartMux(1661) xor i_prn(830)) & (not wbPartMux(1660) xor i_prn(830)) & '1';
    wbMult(2495 downto 2493) := (wbPartMux(1663) xor i_prn(831)) & (not wbPartMux(1662) xor i_prn(831)) & '1';
    wbMult(2498 downto 2496) := (wbPartMux(1665) xor i_prn(832)) & (not wbPartMux(1664) xor i_prn(832)) & '1';
    wbMult(2501 downto 2499) := (wbPartMux(1667) xor i_prn(833)) & (not wbPartMux(1666) xor i_prn(833)) & '1';
    wbMult(2504 downto 2502) := (wbPartMux(1669) xor i_prn(834)) & (not wbPartMux(1668) xor i_prn(834)) & '1';
    wbMult(2507 downto 2505) := (wbPartMux(1671) xor i_prn(835)) & (not wbPartMux(1670) xor i_prn(835)) & '1';
    wbMult(2510 downto 2508) := (wbPartMux(1673) xor i_prn(836)) & (not wbPartMux(1672) xor i_prn(836)) & '1';
    wbMult(2513 downto 2511) := (wbPartMux(1675) xor i_prn(837)) & (not wbPartMux(1674) xor i_prn(837)) & '1';
    wbMult(2516 downto 2514) := (wbPartMux(1677) xor i_prn(838)) & (not wbPartMux(1676) xor i_prn(838)) & '1';
    wbMult(2519 downto 2517) := (wbPartMux(1679) xor i_prn(839)) & (not wbPartMux(1678) xor i_prn(839)) & '1';
    wbMult(2522 downto 2520) := (wbPartMux(1681) xor i_prn(840)) & (not wbPartMux(1680) xor i_prn(840)) & '1';
    wbMult(2525 downto 2523) := (wbPartMux(1683) xor i_prn(841)) & (not wbPartMux(1682) xor i_prn(841)) & '1';
    wbMult(2528 downto 2526) := (wbPartMux(1685) xor i_prn(842)) & (not wbPartMux(1684) xor i_prn(842)) & '1';
    wbMult(2531 downto 2529) := (wbPartMux(1687) xor i_prn(843)) & (not wbPartMux(1686) xor i_prn(843)) & '1';
    wbMult(2534 downto 2532) := (wbPartMux(1689) xor i_prn(844)) & (not wbPartMux(1688) xor i_prn(844)) & '1';
    wbMult(2537 downto 2535) := (wbPartMux(1691) xor i_prn(845)) & (not wbPartMux(1690) xor i_prn(845)) & '1';
    wbMult(2540 downto 2538) := (wbPartMux(1693) xor i_prn(846)) & (not wbPartMux(1692) xor i_prn(846)) & '1';
    wbMult(2543 downto 2541) := (wbPartMux(1695) xor i_prn(847)) & (not wbPartMux(1694) xor i_prn(847)) & '1';
    wbMult(2546 downto 2544) := (wbPartMux(1697) xor i_prn(848)) & (not wbPartMux(1696) xor i_prn(848)) & '1';
    wbMult(2549 downto 2547) := (wbPartMux(1699) xor i_prn(849)) & (not wbPartMux(1698) xor i_prn(849)) & '1';
    wbMult(2552 downto 2550) := (wbPartMux(1701) xor i_prn(850)) & (not wbPartMux(1700) xor i_prn(850)) & '1';
    wbMult(2555 downto 2553) := (wbPartMux(1703) xor i_prn(851)) & (not wbPartMux(1702) xor i_prn(851)) & '1';
    wbMult(2558 downto 2556) := (wbPartMux(1705) xor i_prn(852)) & (not wbPartMux(1704) xor i_prn(852)) & '1';
    wbMult(2561 downto 2559) := (wbPartMux(1707) xor i_prn(853)) & (not wbPartMux(1706) xor i_prn(853)) & '1';
    wbMult(2564 downto 2562) := (wbPartMux(1709) xor i_prn(854)) & (not wbPartMux(1708) xor i_prn(854)) & '1';
    wbMult(2567 downto 2565) := (wbPartMux(1711) xor i_prn(855)) & (not wbPartMux(1710) xor i_prn(855)) & '1';
    wbMult(2570 downto 2568) := (wbPartMux(1713) xor i_prn(856)) & (not wbPartMux(1712) xor i_prn(856)) & '1';
    wbMult(2573 downto 2571) := (wbPartMux(1715) xor i_prn(857)) & (not wbPartMux(1714) xor i_prn(857)) & '1';
    wbMult(2576 downto 2574) := (wbPartMux(1717) xor i_prn(858)) & (not wbPartMux(1716) xor i_prn(858)) & '1';
    wbMult(2579 downto 2577) := (wbPartMux(1719) xor i_prn(859)) & (not wbPartMux(1718) xor i_prn(859)) & '1';
    wbMult(2582 downto 2580) := (wbPartMux(1721) xor i_prn(860)) & (not wbPartMux(1720) xor i_prn(860)) & '1';
    wbMult(2585 downto 2583) := (wbPartMux(1723) xor i_prn(861)) & (not wbPartMux(1722) xor i_prn(861)) & '1';
    wbMult(2588 downto 2586) := (wbPartMux(1725) xor i_prn(862)) & (not wbPartMux(1724) xor i_prn(862)) & '1';
    wbMult(2591 downto 2589) := (wbPartMux(1727) xor i_prn(863)) & (not wbPartMux(1726) xor i_prn(863)) & '1';
    wbMult(2594 downto 2592) := (wbPartMux(1729) xor i_prn(864)) & (not wbPartMux(1728) xor i_prn(864)) & '1';
    wbMult(2597 downto 2595) := (wbPartMux(1731) xor i_prn(865)) & (not wbPartMux(1730) xor i_prn(865)) & '1';
    wbMult(2600 downto 2598) := (wbPartMux(1733) xor i_prn(866)) & (not wbPartMux(1732) xor i_prn(866)) & '1';
    wbMult(2603 downto 2601) := (wbPartMux(1735) xor i_prn(867)) & (not wbPartMux(1734) xor i_prn(867)) & '1';
    wbMult(2606 downto 2604) := (wbPartMux(1737) xor i_prn(868)) & (not wbPartMux(1736) xor i_prn(868)) & '1';
    wbMult(2609 downto 2607) := (wbPartMux(1739) xor i_prn(869)) & (not wbPartMux(1738) xor i_prn(869)) & '1';
    wbMult(2612 downto 2610) := (wbPartMux(1741) xor i_prn(870)) & (not wbPartMux(1740) xor i_prn(870)) & '1';
    wbMult(2615 downto 2613) := (wbPartMux(1743) xor i_prn(871)) & (not wbPartMux(1742) xor i_prn(871)) & '1';
    wbMult(2618 downto 2616) := (wbPartMux(1745) xor i_prn(872)) & (not wbPartMux(1744) xor i_prn(872)) & '1';
    wbMult(2621 downto 2619) := (wbPartMux(1747) xor i_prn(873)) & (not wbPartMux(1746) xor i_prn(873)) & '1';
    wbMult(2624 downto 2622) := (wbPartMux(1749) xor i_prn(874)) & (not wbPartMux(1748) xor i_prn(874)) & '1';
    wbMult(2627 downto 2625) := (wbPartMux(1751) xor i_prn(875)) & (not wbPartMux(1750) xor i_prn(875)) & '1';
    wbMult(2630 downto 2628) := (wbPartMux(1753) xor i_prn(876)) & (not wbPartMux(1752) xor i_prn(876)) & '1';
    wbMult(2633 downto 2631) := (wbPartMux(1755) xor i_prn(877)) & (not wbPartMux(1754) xor i_prn(877)) & '1';
    wbMult(2636 downto 2634) := (wbPartMux(1757) xor i_prn(878)) & (not wbPartMux(1756) xor i_prn(878)) & '1';
    wbMult(2639 downto 2637) := (wbPartMux(1759) xor i_prn(879)) & (not wbPartMux(1758) xor i_prn(879)) & '1';
    wbMult(2642 downto 2640) := (wbPartMux(1761) xor i_prn(880)) & (not wbPartMux(1760) xor i_prn(880)) & '1';
    wbMult(2645 downto 2643) := (wbPartMux(1763) xor i_prn(881)) & (not wbPartMux(1762) xor i_prn(881)) & '1';
    wbMult(2648 downto 2646) := (wbPartMux(1765) xor i_prn(882)) & (not wbPartMux(1764) xor i_prn(882)) & '1';
    wbMult(2651 downto 2649) := (wbPartMux(1767) xor i_prn(883)) & (not wbPartMux(1766) xor i_prn(883)) & '1';
    wbMult(2654 downto 2652) := (wbPartMux(1769) xor i_prn(884)) & (not wbPartMux(1768) xor i_prn(884)) & '1';
    wbMult(2657 downto 2655) := (wbPartMux(1771) xor i_prn(885)) & (not wbPartMux(1770) xor i_prn(885)) & '1';
    wbMult(2660 downto 2658) := (wbPartMux(1773) xor i_prn(886)) & (not wbPartMux(1772) xor i_prn(886)) & '1';
    wbMult(2663 downto 2661) := (wbPartMux(1775) xor i_prn(887)) & (not wbPartMux(1774) xor i_prn(887)) & '1';
    wbMult(2666 downto 2664) := (wbPartMux(1777) xor i_prn(888)) & (not wbPartMux(1776) xor i_prn(888)) & '1';
    wbMult(2669 downto 2667) := (wbPartMux(1779) xor i_prn(889)) & (not wbPartMux(1778) xor i_prn(889)) & '1';
    wbMult(2672 downto 2670) := (wbPartMux(1781) xor i_prn(890)) & (not wbPartMux(1780) xor i_prn(890)) & '1';
    wbMult(2675 downto 2673) := (wbPartMux(1783) xor i_prn(891)) & (not wbPartMux(1782) xor i_prn(891)) & '1';
    wbMult(2678 downto 2676) := (wbPartMux(1785) xor i_prn(892)) & (not wbPartMux(1784) xor i_prn(892)) & '1';
    wbMult(2681 downto 2679) := (wbPartMux(1787) xor i_prn(893)) & (not wbPartMux(1786) xor i_prn(893)) & '1';
    wbMult(2684 downto 2682) := (wbPartMux(1789) xor i_prn(894)) & (not wbPartMux(1788) xor i_prn(894)) & '1';
    wbMult(2687 downto 2685) := (wbPartMux(1791) xor i_prn(895)) & (not wbPartMux(1790) xor i_prn(895)) & '1';
    wbMult(2690 downto 2688) := (wbPartMux(1793) xor i_prn(896)) & (not wbPartMux(1792) xor i_prn(896)) & '1';
    wbMult(2693 downto 2691) := (wbPartMux(1795) xor i_prn(897)) & (not wbPartMux(1794) xor i_prn(897)) & '1';
    wbMult(2696 downto 2694) := (wbPartMux(1797) xor i_prn(898)) & (not wbPartMux(1796) xor i_prn(898)) & '1';
    wbMult(2699 downto 2697) := (wbPartMux(1799) xor i_prn(899)) & (not wbPartMux(1798) xor i_prn(899)) & '1';
    wbMult(2702 downto 2700) := (wbPartMux(1801) xor i_prn(900)) & (not wbPartMux(1800) xor i_prn(900)) & '1';
    wbMult(2705 downto 2703) := (wbPartMux(1803) xor i_prn(901)) & (not wbPartMux(1802) xor i_prn(901)) & '1';
    wbMult(2708 downto 2706) := (wbPartMux(1805) xor i_prn(902)) & (not wbPartMux(1804) xor i_prn(902)) & '1';
    wbMult(2711 downto 2709) := (wbPartMux(1807) xor i_prn(903)) & (not wbPartMux(1806) xor i_prn(903)) & '1';
    wbMult(2714 downto 2712) := (wbPartMux(1809) xor i_prn(904)) & (not wbPartMux(1808) xor i_prn(904)) & '1';
    wbMult(2717 downto 2715) := (wbPartMux(1811) xor i_prn(905)) & (not wbPartMux(1810) xor i_prn(905)) & '1';
    wbMult(2720 downto 2718) := (wbPartMux(1813) xor i_prn(906)) & (not wbPartMux(1812) xor i_prn(906)) & '1';
    wbMult(2723 downto 2721) := (wbPartMux(1815) xor i_prn(907)) & (not wbPartMux(1814) xor i_prn(907)) & '1';
    wbMult(2726 downto 2724) := (wbPartMux(1817) xor i_prn(908)) & (not wbPartMux(1816) xor i_prn(908)) & '1';
    wbMult(2729 downto 2727) := (wbPartMux(1819) xor i_prn(909)) & (not wbPartMux(1818) xor i_prn(909)) & '1';
    wbMult(2732 downto 2730) := (wbPartMux(1821) xor i_prn(910)) & (not wbPartMux(1820) xor i_prn(910)) & '1';
    wbMult(2735 downto 2733) := (wbPartMux(1823) xor i_prn(911)) & (not wbPartMux(1822) xor i_prn(911)) & '1';
    wbMult(2738 downto 2736) := (wbPartMux(1825) xor i_prn(912)) & (not wbPartMux(1824) xor i_prn(912)) & '1';
    wbMult(2741 downto 2739) := (wbPartMux(1827) xor i_prn(913)) & (not wbPartMux(1826) xor i_prn(913)) & '1';
    wbMult(2744 downto 2742) := (wbPartMux(1829) xor i_prn(914)) & (not wbPartMux(1828) xor i_prn(914)) & '1';
    wbMult(2747 downto 2745) := (wbPartMux(1831) xor i_prn(915)) & (not wbPartMux(1830) xor i_prn(915)) & '1';
    wbMult(2750 downto 2748) := (wbPartMux(1833) xor i_prn(916)) & (not wbPartMux(1832) xor i_prn(916)) & '1';
    wbMult(2753 downto 2751) := (wbPartMux(1835) xor i_prn(917)) & (not wbPartMux(1834) xor i_prn(917)) & '1';
    wbMult(2756 downto 2754) := (wbPartMux(1837) xor i_prn(918)) & (not wbPartMux(1836) xor i_prn(918)) & '1';
    wbMult(2759 downto 2757) := (wbPartMux(1839) xor i_prn(919)) & (not wbPartMux(1838) xor i_prn(919)) & '1';
    wbMult(2762 downto 2760) := (wbPartMux(1841) xor i_prn(920)) & (not wbPartMux(1840) xor i_prn(920)) & '1';
    wbMult(2765 downto 2763) := (wbPartMux(1843) xor i_prn(921)) & (not wbPartMux(1842) xor i_prn(921)) & '1';
    wbMult(2768 downto 2766) := (wbPartMux(1845) xor i_prn(922)) & (not wbPartMux(1844) xor i_prn(922)) & '1';
    wbMult(2771 downto 2769) := (wbPartMux(1847) xor i_prn(923)) & (not wbPartMux(1846) xor i_prn(923)) & '1';
    wbMult(2774 downto 2772) := (wbPartMux(1849) xor i_prn(924)) & (not wbPartMux(1848) xor i_prn(924)) & '1';
    wbMult(2777 downto 2775) := (wbPartMux(1851) xor i_prn(925)) & (not wbPartMux(1850) xor i_prn(925)) & '1';
    wbMult(2780 downto 2778) := (wbPartMux(1853) xor i_prn(926)) & (not wbPartMux(1852) xor i_prn(926)) & '1';
    wbMult(2783 downto 2781) := (wbPartMux(1855) xor i_prn(927)) & (not wbPartMux(1854) xor i_prn(927)) & '1';
    wbMult(2786 downto 2784) := (wbPartMux(1857) xor i_prn(928)) & (not wbPartMux(1856) xor i_prn(928)) & '1';
    wbMult(2789 downto 2787) := (wbPartMux(1859) xor i_prn(929)) & (not wbPartMux(1858) xor i_prn(929)) & '1';
    wbMult(2792 downto 2790) := (wbPartMux(1861) xor i_prn(930)) & (not wbPartMux(1860) xor i_prn(930)) & '1';
    wbMult(2795 downto 2793) := (wbPartMux(1863) xor i_prn(931)) & (not wbPartMux(1862) xor i_prn(931)) & '1';
    wbMult(2798 downto 2796) := (wbPartMux(1865) xor i_prn(932)) & (not wbPartMux(1864) xor i_prn(932)) & '1';
    wbMult(2801 downto 2799) := (wbPartMux(1867) xor i_prn(933)) & (not wbPartMux(1866) xor i_prn(933)) & '1';
    wbMult(2804 downto 2802) := (wbPartMux(1869) xor i_prn(934)) & (not wbPartMux(1868) xor i_prn(934)) & '1';
    wbMult(2807 downto 2805) := (wbPartMux(1871) xor i_prn(935)) & (not wbPartMux(1870) xor i_prn(935)) & '1';
    wbMult(2810 downto 2808) := (wbPartMux(1873) xor i_prn(936)) & (not wbPartMux(1872) xor i_prn(936)) & '1';
    wbMult(2813 downto 2811) := (wbPartMux(1875) xor i_prn(937)) & (not wbPartMux(1874) xor i_prn(937)) & '1';
    wbMult(2816 downto 2814) := (wbPartMux(1877) xor i_prn(938)) & (not wbPartMux(1876) xor i_prn(938)) & '1';
    wbMult(2819 downto 2817) := (wbPartMux(1879) xor i_prn(939)) & (not wbPartMux(1878) xor i_prn(939)) & '1';
    wbMult(2822 downto 2820) := (wbPartMux(1881) xor i_prn(940)) & (not wbPartMux(1880) xor i_prn(940)) & '1';
    wbMult(2825 downto 2823) := (wbPartMux(1883) xor i_prn(941)) & (not wbPartMux(1882) xor i_prn(941)) & '1';
    wbMult(2828 downto 2826) := (wbPartMux(1885) xor i_prn(942)) & (not wbPartMux(1884) xor i_prn(942)) & '1';
    wbMult(2831 downto 2829) := (wbPartMux(1887) xor i_prn(943)) & (not wbPartMux(1886) xor i_prn(943)) & '1';
    wbMult(2834 downto 2832) := (wbPartMux(1889) xor i_prn(944)) & (not wbPartMux(1888) xor i_prn(944)) & '1';
    wbMult(2837 downto 2835) := (wbPartMux(1891) xor i_prn(945)) & (not wbPartMux(1890) xor i_prn(945)) & '1';
    wbMult(2840 downto 2838) := (wbPartMux(1893) xor i_prn(946)) & (not wbPartMux(1892) xor i_prn(946)) & '1';
    wbMult(2843 downto 2841) := (wbPartMux(1895) xor i_prn(947)) & (not wbPartMux(1894) xor i_prn(947)) & '1';
    wbMult(2846 downto 2844) := (wbPartMux(1897) xor i_prn(948)) & (not wbPartMux(1896) xor i_prn(948)) & '1';
    wbMult(2849 downto 2847) := (wbPartMux(1899) xor i_prn(949)) & (not wbPartMux(1898) xor i_prn(949)) & '1';
    wbMult(2852 downto 2850) := (wbPartMux(1901) xor i_prn(950)) & (not wbPartMux(1900) xor i_prn(950)) & '1';
    wbMult(2855 downto 2853) := (wbPartMux(1903) xor i_prn(951)) & (not wbPartMux(1902) xor i_prn(951)) & '1';
    wbMult(2858 downto 2856) := (wbPartMux(1905) xor i_prn(952)) & (not wbPartMux(1904) xor i_prn(952)) & '1';
    wbMult(2861 downto 2859) := (wbPartMux(1907) xor i_prn(953)) & (not wbPartMux(1906) xor i_prn(953)) & '1';
    wbMult(2864 downto 2862) := (wbPartMux(1909) xor i_prn(954)) & (not wbPartMux(1908) xor i_prn(954)) & '1';
    wbMult(2867 downto 2865) := (wbPartMux(1911) xor i_prn(955)) & (not wbPartMux(1910) xor i_prn(955)) & '1';
    wbMult(2870 downto 2868) := (wbPartMux(1913) xor i_prn(956)) & (not wbPartMux(1912) xor i_prn(956)) & '1';
    wbMult(2873 downto 2871) := (wbPartMux(1915) xor i_prn(957)) & (not wbPartMux(1914) xor i_prn(957)) & '1';
    wbMult(2876 downto 2874) := (wbPartMux(1917) xor i_prn(958)) & (not wbPartMux(1916) xor i_prn(958)) & '1';
    wbMult(2879 downto 2877) := (wbPartMux(1919) xor i_prn(959)) & (not wbPartMux(1918) xor i_prn(959)) & '1';
    wbMult(2882 downto 2880) := (wbPartMux(1921) xor i_prn(960)) & (not wbPartMux(1920) xor i_prn(960)) & '1';
    wbMult(2885 downto 2883) := (wbPartMux(1923) xor i_prn(961)) & (not wbPartMux(1922) xor i_prn(961)) & '1';
    wbMult(2888 downto 2886) := (wbPartMux(1925) xor i_prn(962)) & (not wbPartMux(1924) xor i_prn(962)) & '1';
    wbMult(2891 downto 2889) := (wbPartMux(1927) xor i_prn(963)) & (not wbPartMux(1926) xor i_prn(963)) & '1';
    wbMult(2894 downto 2892) := (wbPartMux(1929) xor i_prn(964)) & (not wbPartMux(1928) xor i_prn(964)) & '1';
    wbMult(2897 downto 2895) := (wbPartMux(1931) xor i_prn(965)) & (not wbPartMux(1930) xor i_prn(965)) & '1';
    wbMult(2900 downto 2898) := (wbPartMux(1933) xor i_prn(966)) & (not wbPartMux(1932) xor i_prn(966)) & '1';
    wbMult(2903 downto 2901) := (wbPartMux(1935) xor i_prn(967)) & (not wbPartMux(1934) xor i_prn(967)) & '1';
    wbMult(2906 downto 2904) := (wbPartMux(1937) xor i_prn(968)) & (not wbPartMux(1936) xor i_prn(968)) & '1';
    wbMult(2909 downto 2907) := (wbPartMux(1939) xor i_prn(969)) & (not wbPartMux(1938) xor i_prn(969)) & '1';
    wbMult(2912 downto 2910) := (wbPartMux(1941) xor i_prn(970)) & (not wbPartMux(1940) xor i_prn(970)) & '1';
    wbMult(2915 downto 2913) := (wbPartMux(1943) xor i_prn(971)) & (not wbPartMux(1942) xor i_prn(971)) & '1';
    wbMult(2918 downto 2916) := (wbPartMux(1945) xor i_prn(972)) & (not wbPartMux(1944) xor i_prn(972)) & '1';
    wbMult(2921 downto 2919) := (wbPartMux(1947) xor i_prn(973)) & (not wbPartMux(1946) xor i_prn(973)) & '1';
    wbMult(2924 downto 2922) := (wbPartMux(1949) xor i_prn(974)) & (not wbPartMux(1948) xor i_prn(974)) & '1';
    wbMult(2927 downto 2925) := (wbPartMux(1951) xor i_prn(975)) & (not wbPartMux(1950) xor i_prn(975)) & '1';
    wbMult(2930 downto 2928) := (wbPartMux(1953) xor i_prn(976)) & (not wbPartMux(1952) xor i_prn(976)) & '1';
    wbMult(2933 downto 2931) := (wbPartMux(1955) xor i_prn(977)) & (not wbPartMux(1954) xor i_prn(977)) & '1';
    wbMult(2936 downto 2934) := (wbPartMux(1957) xor i_prn(978)) & (not wbPartMux(1956) xor i_prn(978)) & '1';
    wbMult(2939 downto 2937) := (wbPartMux(1959) xor i_prn(979)) & (not wbPartMux(1958) xor i_prn(979)) & '1';
    wbMult(2942 downto 2940) := (wbPartMux(1961) xor i_prn(980)) & (not wbPartMux(1960) xor i_prn(980)) & '1';
    wbMult(2945 downto 2943) := (wbPartMux(1963) xor i_prn(981)) & (not wbPartMux(1962) xor i_prn(981)) & '1';
    wbMult(2948 downto 2946) := (wbPartMux(1965) xor i_prn(982)) & (not wbPartMux(1964) xor i_prn(982)) & '1';
    wbMult(2951 downto 2949) := (wbPartMux(1967) xor i_prn(983)) & (not wbPartMux(1966) xor i_prn(983)) & '1';
    wbMult(2954 downto 2952) := (wbPartMux(1969) xor i_prn(984)) & (not wbPartMux(1968) xor i_prn(984)) & '1';
    wbMult(2957 downto 2955) := (wbPartMux(1971) xor i_prn(985)) & (not wbPartMux(1970) xor i_prn(985)) & '1';
    wbMult(2960 downto 2958) := (wbPartMux(1973) xor i_prn(986)) & (not wbPartMux(1972) xor i_prn(986)) & '1';
    wbMult(2963 downto 2961) := (wbPartMux(1975) xor i_prn(987)) & (not wbPartMux(1974) xor i_prn(987)) & '1';
    wbMult(2966 downto 2964) := (wbPartMux(1977) xor i_prn(988)) & (not wbPartMux(1976) xor i_prn(988)) & '1';
    wbMult(2969 downto 2967) := (wbPartMux(1979) xor i_prn(989)) & (not wbPartMux(1978) xor i_prn(989)) & '1';
    wbMult(2972 downto 2970) := (wbPartMux(1981) xor i_prn(990)) & (not wbPartMux(1980) xor i_prn(990)) & '1';
    wbMult(2975 downto 2973) := (wbPartMux(1983) xor i_prn(991)) & (not wbPartMux(1982) xor i_prn(991)) & '1';
    wbMult(2978 downto 2976) := (wbPartMux(1985) xor i_prn(992)) & (not wbPartMux(1984) xor i_prn(992)) & '1';
    wbMult(2981 downto 2979) := (wbPartMux(1987) xor i_prn(993)) & (not wbPartMux(1986) xor i_prn(993)) & '1';
    wbMult(2984 downto 2982) := (wbPartMux(1989) xor i_prn(994)) & (not wbPartMux(1988) xor i_prn(994)) & '1';
    wbMult(2987 downto 2985) := (wbPartMux(1991) xor i_prn(995)) & (not wbPartMux(1990) xor i_prn(995)) & '1';
    wbMult(2990 downto 2988) := (wbPartMux(1993) xor i_prn(996)) & (not wbPartMux(1992) xor i_prn(996)) & '1';
    wbMult(2993 downto 2991) := (wbPartMux(1995) xor i_prn(997)) & (not wbPartMux(1994) xor i_prn(997)) & '1';
    wbMult(2996 downto 2994) := (wbPartMux(1997) xor i_prn(998)) & (not wbPartMux(1996) xor i_prn(998)) & '1';
    wbMult(2999 downto 2997) := (wbPartMux(1999) xor i_prn(999)) & (not wbPartMux(1998) xor i_prn(999)) & '1';
    wbMult(3002 downto 3000) := (wbPartMux(2001) xor i_prn(1000)) & (not wbPartMux(2000) xor i_prn(1000)) & '1';
    wbMult(3005 downto 3003) := (wbPartMux(2003) xor i_prn(1001)) & (not wbPartMux(2002) xor i_prn(1001)) & '1';
    wbMult(3008 downto 3006) := (wbPartMux(2005) xor i_prn(1002)) & (not wbPartMux(2004) xor i_prn(1002)) & '1';
    wbMult(3011 downto 3009) := (wbPartMux(2007) xor i_prn(1003)) & (not wbPartMux(2006) xor i_prn(1003)) & '1';
    wbMult(3014 downto 3012) := (wbPartMux(2009) xor i_prn(1004)) & (not wbPartMux(2008) xor i_prn(1004)) & '1';
    wbMult(3017 downto 3015) := (wbPartMux(2011) xor i_prn(1005)) & (not wbPartMux(2010) xor i_prn(1005)) & '1';
    wbMult(3020 downto 3018) := (wbPartMux(2013) xor i_prn(1006)) & (not wbPartMux(2012) xor i_prn(1006)) & '1';
    wbMult(3023 downto 3021) := (wbPartMux(2015) xor i_prn(1007)) & (not wbPartMux(2014) xor i_prn(1007)) & '1';
    wbMult(3026 downto 3024) := (wbPartMux(2017) xor i_prn(1008)) & (not wbPartMux(2016) xor i_prn(1008)) & '1';
    wbMult(3029 downto 3027) := (wbPartMux(2019) xor i_prn(1009)) & (not wbPartMux(2018) xor i_prn(1009)) & '1';
    wbMult(3032 downto 3030) := (wbPartMux(2021) xor i_prn(1010)) & (not wbPartMux(2020) xor i_prn(1010)) & '1';
    wbMult(3035 downto 3033) := (wbPartMux(2023) xor i_prn(1011)) & (not wbPartMux(2022) xor i_prn(1011)) & '1';
    wbMult(3038 downto 3036) := (wbPartMux(2025) xor i_prn(1012)) & (not wbPartMux(2024) xor i_prn(1012)) & '1';
    wbMult(3041 downto 3039) := (wbPartMux(2027) xor i_prn(1013)) & (not wbPartMux(2026) xor i_prn(1013)) & '1';
    wbMult(3044 downto 3042) := (wbPartMux(2029) xor i_prn(1014)) & (not wbPartMux(2028) xor i_prn(1014)) & '1';
    wbMult(3047 downto 3045) := (wbPartMux(2031) xor i_prn(1015)) & (not wbPartMux(2030) xor i_prn(1015)) & '1';
    wbMult(3050 downto 3048) := (wbPartMux(2033) xor i_prn(1016)) & (not wbPartMux(2032) xor i_prn(1016)) & '1';
    wbMult(3053 downto 3051) := (wbPartMux(2035) xor i_prn(1017)) & (not wbPartMux(2034) xor i_prn(1017)) & '1';
    wbMult(3056 downto 3054) := (wbPartMux(2037) xor i_prn(1018)) & (not wbPartMux(2036) xor i_prn(1018)) & '1';
    wbMult(3059 downto 3057) := (wbPartMux(2039) xor i_prn(1019)) & (not wbPartMux(2038) xor i_prn(1019)) & '1';
    wbMult(3062 downto 3060) := (wbPartMux(2041) xor i_prn(1020)) & (not wbPartMux(2040) xor i_prn(1020)) & '1';
    wbMult(3065 downto 3063) := (wbPartMux(2043) xor i_prn(1021)) & (not wbPartMux(2042) xor i_prn(1021)) & '1';
    wbMult(3068 downto 3066) := (wbPartMux(2045) xor i_prn(1022)) & (not wbPartMux(2044) xor i_prn(1022)) & '1';
    wbMult(3071 downto 3069) := (wbPartMux(2047) xor i_prn(1023)) & (not wbPartMux(2046) xor i_prn(1023)) & '1';


    --if i.ena = '1' then
      v.Lvl1(3 downto 0) := (wbMult(2) & wbMult(2 downto 0)) + (wbMult(5) & wbMult(5 downto 3));
      v.Lvl1(7 downto 4) := (wbMult(8) & wbMult(8 downto 6)) + (wbMult(11) & wbMult(11 downto 9));
      v.Lvl1(11 downto 8) := (wbMult(14) & wbMult(14 downto 12)) + (wbMult(17) & wbMult(17 downto 15));
      v.Lvl1(15 downto 12) := (wbMult(20) & wbMult(20 downto 18)) + (wbMult(23) & wbMult(23 downto 21));
      v.Lvl1(19 downto 16) := (wbMult(26) & wbMult(26 downto 24)) + (wbMult(29) & wbMult(29 downto 27));
      v.Lvl1(23 downto 20) := (wbMult(32) & wbMult(32 downto 30)) + (wbMult(35) & wbMult(35 downto 33));
      v.Lvl1(27 downto 24) := (wbMult(38) & wbMult(38 downto 36)) + (wbMult(41) & wbMult(41 downto 39));
      v.Lvl1(31 downto 28) := (wbMult(44) & wbMult(44 downto 42)) + (wbMult(47) & wbMult(47 downto 45));
      v.Lvl1(35 downto 32) := (wbMult(50) & wbMult(50 downto 48)) + (wbMult(53) & wbMult(53 downto 51));
      v.Lvl1(39 downto 36) := (wbMult(56) & wbMult(56 downto 54)) + (wbMult(59) & wbMult(59 downto 57));
      v.Lvl1(43 downto 40) := (wbMult(62) & wbMult(62 downto 60)) + (wbMult(65) & wbMult(65 downto 63));
      v.Lvl1(47 downto 44) := (wbMult(68) & wbMult(68 downto 66)) + (wbMult(71) & wbMult(71 downto 69));
      v.Lvl1(51 downto 48) := (wbMult(74) & wbMult(74 downto 72)) + (wbMult(77) & wbMult(77 downto 75));
      v.Lvl1(55 downto 52) := (wbMult(80) & wbMult(80 downto 78)) + (wbMult(83) & wbMult(83 downto 81));
      v.Lvl1(59 downto 56) := (wbMult(86) & wbMult(86 downto 84)) + (wbMult(89) & wbMult(89 downto 87));
      v.Lvl1(63 downto 60) := (wbMult(92) & wbMult(92 downto 90)) + (wbMult(95) & wbMult(95 downto 93));
      v.Lvl1(67 downto 64) := (wbMult(98) & wbMult(98 downto 96)) + (wbMult(101) & wbMult(101 downto 99));
      v.Lvl1(71 downto 68) := (wbMult(104) & wbMult(104 downto 102)) + (wbMult(107) & wbMult(107 downto 105));
      v.Lvl1(75 downto 72) := (wbMult(110) & wbMult(110 downto 108)) + (wbMult(113) & wbMult(113 downto 111));
      v.Lvl1(79 downto 76) := (wbMult(116) & wbMult(116 downto 114)) + (wbMult(119) & wbMult(119 downto 117));
      v.Lvl1(83 downto 80) := (wbMult(122) & wbMult(122 downto 120)) + (wbMult(125) & wbMult(125 downto 123));
      v.Lvl1(87 downto 84) := (wbMult(128) & wbMult(128 downto 126)) + (wbMult(131) & wbMult(131 downto 129));
      v.Lvl1(91 downto 88) := (wbMult(134) & wbMult(134 downto 132)) + (wbMult(137) & wbMult(137 downto 135));
      v.Lvl1(95 downto 92) := (wbMult(140) & wbMult(140 downto 138)) + (wbMult(143) & wbMult(143 downto 141));
      v.Lvl1(99 downto 96) := (wbMult(146) & wbMult(146 downto 144)) + (wbMult(149) & wbMult(149 downto 147));
      v.Lvl1(103 downto 100) := (wbMult(152) & wbMult(152 downto 150)) + (wbMult(155) & wbMult(155 downto 153));
      v.Lvl1(107 downto 104) := (wbMult(158) & wbMult(158 downto 156)) + (wbMult(161) & wbMult(161 downto 159));
      v.Lvl1(111 downto 108) := (wbMult(164) & wbMult(164 downto 162)) + (wbMult(167) & wbMult(167 downto 165));
      v.Lvl1(115 downto 112) := (wbMult(170) & wbMult(170 downto 168)) + (wbMult(173) & wbMult(173 downto 171));
      v.Lvl1(119 downto 116) := (wbMult(176) & wbMult(176 downto 174)) + (wbMult(179) & wbMult(179 downto 177));
      v.Lvl1(123 downto 120) := (wbMult(182) & wbMult(182 downto 180)) + (wbMult(185) & wbMult(185 downto 183));
      v.Lvl1(127 downto 124) := (wbMult(188) & wbMult(188 downto 186)) + (wbMult(191) & wbMult(191 downto 189));
      v.Lvl1(131 downto 128) := (wbMult(194) & wbMult(194 downto 192)) + (wbMult(197) & wbMult(197 downto 195));
      v.Lvl1(135 downto 132) := (wbMult(200) & wbMult(200 downto 198)) + (wbMult(203) & wbMult(203 downto 201));
      v.Lvl1(139 downto 136) := (wbMult(206) & wbMult(206 downto 204)) + (wbMult(209) & wbMult(209 downto 207));
      v.Lvl1(143 downto 140) := (wbMult(212) & wbMult(212 downto 210)) + (wbMult(215) & wbMult(215 downto 213));
      v.Lvl1(147 downto 144) := (wbMult(218) & wbMult(218 downto 216)) + (wbMult(221) & wbMult(221 downto 219));
      v.Lvl1(151 downto 148) := (wbMult(224) & wbMult(224 downto 222)) + (wbMult(227) & wbMult(227 downto 225));
      v.Lvl1(155 downto 152) := (wbMult(230) & wbMult(230 downto 228)) + (wbMult(233) & wbMult(233 downto 231));
      v.Lvl1(159 downto 156) := (wbMult(236) & wbMult(236 downto 234)) + (wbMult(239) & wbMult(239 downto 237));
      v.Lvl1(163 downto 160) := (wbMult(242) & wbMult(242 downto 240)) + (wbMult(245) & wbMult(245 downto 243));
      v.Lvl1(167 downto 164) := (wbMult(248) & wbMult(248 downto 246)) + (wbMult(251) & wbMult(251 downto 249));
      v.Lvl1(171 downto 168) := (wbMult(254) & wbMult(254 downto 252)) + (wbMult(257) & wbMult(257 downto 255));
      v.Lvl1(175 downto 172) := (wbMult(260) & wbMult(260 downto 258)) + (wbMult(263) & wbMult(263 downto 261));
      v.Lvl1(179 downto 176) := (wbMult(266) & wbMult(266 downto 264)) + (wbMult(269) & wbMult(269 downto 267));
      v.Lvl1(183 downto 180) := (wbMult(272) & wbMult(272 downto 270)) + (wbMult(275) & wbMult(275 downto 273));
      v.Lvl1(187 downto 184) := (wbMult(278) & wbMult(278 downto 276)) + (wbMult(281) & wbMult(281 downto 279));
      v.Lvl1(191 downto 188) := (wbMult(284) & wbMult(284 downto 282)) + (wbMult(287) & wbMult(287 downto 285));
      v.Lvl1(195 downto 192) := (wbMult(290) & wbMult(290 downto 288)) + (wbMult(293) & wbMult(293 downto 291));
      v.Lvl1(199 downto 196) := (wbMult(296) & wbMult(296 downto 294)) + (wbMult(299) & wbMult(299 downto 297));
      v.Lvl1(203 downto 200) := (wbMult(302) & wbMult(302 downto 300)) + (wbMult(305) & wbMult(305 downto 303));
      v.Lvl1(207 downto 204) := (wbMult(308) & wbMult(308 downto 306)) + (wbMult(311) & wbMult(311 downto 309));
      v.Lvl1(211 downto 208) := (wbMult(314) & wbMult(314 downto 312)) + (wbMult(317) & wbMult(317 downto 315));
      v.Lvl1(215 downto 212) := (wbMult(320) & wbMult(320 downto 318)) + (wbMult(323) & wbMult(323 downto 321));
      v.Lvl1(219 downto 216) := (wbMult(326) & wbMult(326 downto 324)) + (wbMult(329) & wbMult(329 downto 327));
      v.Lvl1(223 downto 220) := (wbMult(332) & wbMult(332 downto 330)) + (wbMult(335) & wbMult(335 downto 333));
      v.Lvl1(227 downto 224) := (wbMult(338) & wbMult(338 downto 336)) + (wbMult(341) & wbMult(341 downto 339));
      v.Lvl1(231 downto 228) := (wbMult(344) & wbMult(344 downto 342)) + (wbMult(347) & wbMult(347 downto 345));
      v.Lvl1(235 downto 232) := (wbMult(350) & wbMult(350 downto 348)) + (wbMult(353) & wbMult(353 downto 351));
      v.Lvl1(239 downto 236) := (wbMult(356) & wbMult(356 downto 354)) + (wbMult(359) & wbMult(359 downto 357));
      v.Lvl1(243 downto 240) := (wbMult(362) & wbMult(362 downto 360)) + (wbMult(365) & wbMult(365 downto 363));
      v.Lvl1(247 downto 244) := (wbMult(368) & wbMult(368 downto 366)) + (wbMult(371) & wbMult(371 downto 369));
      v.Lvl1(251 downto 248) := (wbMult(374) & wbMult(374 downto 372)) + (wbMult(377) & wbMult(377 downto 375));
      v.Lvl1(255 downto 252) := (wbMult(380) & wbMult(380 downto 378)) + (wbMult(383) & wbMult(383 downto 381));
      v.Lvl1(259 downto 256) := (wbMult(386) & wbMult(386 downto 384)) + (wbMult(389) & wbMult(389 downto 387));
      v.Lvl1(263 downto 260) := (wbMult(392) & wbMult(392 downto 390)) + (wbMult(395) & wbMult(395 downto 393));
      v.Lvl1(267 downto 264) := (wbMult(398) & wbMult(398 downto 396)) + (wbMult(401) & wbMult(401 downto 399));
      v.Lvl1(271 downto 268) := (wbMult(404) & wbMult(404 downto 402)) + (wbMult(407) & wbMult(407 downto 405));
      v.Lvl1(275 downto 272) := (wbMult(410) & wbMult(410 downto 408)) + (wbMult(413) & wbMult(413 downto 411));
      v.Lvl1(279 downto 276) := (wbMult(416) & wbMult(416 downto 414)) + (wbMult(419) & wbMult(419 downto 417));
      v.Lvl1(283 downto 280) := (wbMult(422) & wbMult(422 downto 420)) + (wbMult(425) & wbMult(425 downto 423));
      v.Lvl1(287 downto 284) := (wbMult(428) & wbMult(428 downto 426)) + (wbMult(431) & wbMult(431 downto 429));
      v.Lvl1(291 downto 288) := (wbMult(434) & wbMult(434 downto 432)) + (wbMult(437) & wbMult(437 downto 435));
      v.Lvl1(295 downto 292) := (wbMult(440) & wbMult(440 downto 438)) + (wbMult(443) & wbMult(443 downto 441));
      v.Lvl1(299 downto 296) := (wbMult(446) & wbMult(446 downto 444)) + (wbMult(449) & wbMult(449 downto 447));
      v.Lvl1(303 downto 300) := (wbMult(452) & wbMult(452 downto 450)) + (wbMult(455) & wbMult(455 downto 453));
      v.Lvl1(307 downto 304) := (wbMult(458) & wbMult(458 downto 456)) + (wbMult(461) & wbMult(461 downto 459));
      v.Lvl1(311 downto 308) := (wbMult(464) & wbMult(464 downto 462)) + (wbMult(467) & wbMult(467 downto 465));
      v.Lvl1(315 downto 312) := (wbMult(470) & wbMult(470 downto 468)) + (wbMult(473) & wbMult(473 downto 471));
      v.Lvl1(319 downto 316) := (wbMult(476) & wbMult(476 downto 474)) + (wbMult(479) & wbMult(479 downto 477));
      v.Lvl1(323 downto 320) := (wbMult(482) & wbMult(482 downto 480)) + (wbMult(485) & wbMult(485 downto 483));
      v.Lvl1(327 downto 324) := (wbMult(488) & wbMult(488 downto 486)) + (wbMult(491) & wbMult(491 downto 489));
      v.Lvl1(331 downto 328) := (wbMult(494) & wbMult(494 downto 492)) + (wbMult(497) & wbMult(497 downto 495));
      v.Lvl1(335 downto 332) := (wbMult(500) & wbMult(500 downto 498)) + (wbMult(503) & wbMult(503 downto 501));
      v.Lvl1(339 downto 336) := (wbMult(506) & wbMult(506 downto 504)) + (wbMult(509) & wbMult(509 downto 507));
      v.Lvl1(343 downto 340) := (wbMult(512) & wbMult(512 downto 510)) + (wbMult(515) & wbMult(515 downto 513));
      v.Lvl1(347 downto 344) := (wbMult(518) & wbMult(518 downto 516)) + (wbMult(521) & wbMult(521 downto 519));
      v.Lvl1(351 downto 348) := (wbMult(524) & wbMult(524 downto 522)) + (wbMult(527) & wbMult(527 downto 525));
      v.Lvl1(355 downto 352) := (wbMult(530) & wbMult(530 downto 528)) + (wbMult(533) & wbMult(533 downto 531));
      v.Lvl1(359 downto 356) := (wbMult(536) & wbMult(536 downto 534)) + (wbMult(539) & wbMult(539 downto 537));
      v.Lvl1(363 downto 360) := (wbMult(542) & wbMult(542 downto 540)) + (wbMult(545) & wbMult(545 downto 543));
      v.Lvl1(367 downto 364) := (wbMult(548) & wbMult(548 downto 546)) + (wbMult(551) & wbMult(551 downto 549));
      v.Lvl1(371 downto 368) := (wbMult(554) & wbMult(554 downto 552)) + (wbMult(557) & wbMult(557 downto 555));
      v.Lvl1(375 downto 372) := (wbMult(560) & wbMult(560 downto 558)) + (wbMult(563) & wbMult(563 downto 561));
      v.Lvl1(379 downto 376) := (wbMult(566) & wbMult(566 downto 564)) + (wbMult(569) & wbMult(569 downto 567));
      v.Lvl1(383 downto 380) := (wbMult(572) & wbMult(572 downto 570)) + (wbMult(575) & wbMult(575 downto 573));
      v.Lvl1(387 downto 384) := (wbMult(578) & wbMult(578 downto 576)) + (wbMult(581) & wbMult(581 downto 579));
      v.Lvl1(391 downto 388) := (wbMult(584) & wbMult(584 downto 582)) + (wbMult(587) & wbMult(587 downto 585));
      v.Lvl1(395 downto 392) := (wbMult(590) & wbMult(590 downto 588)) + (wbMult(593) & wbMult(593 downto 591));
      v.Lvl1(399 downto 396) := (wbMult(596) & wbMult(596 downto 594)) + (wbMult(599) & wbMult(599 downto 597));
      v.Lvl1(403 downto 400) := (wbMult(602) & wbMult(602 downto 600)) + (wbMult(605) & wbMult(605 downto 603));
      v.Lvl1(407 downto 404) := (wbMult(608) & wbMult(608 downto 606)) + (wbMult(611) & wbMult(611 downto 609));
      v.Lvl1(411 downto 408) := (wbMult(614) & wbMult(614 downto 612)) + (wbMult(617) & wbMult(617 downto 615));
      v.Lvl1(415 downto 412) := (wbMult(620) & wbMult(620 downto 618)) + (wbMult(623) & wbMult(623 downto 621));
      v.Lvl1(419 downto 416) := (wbMult(626) & wbMult(626 downto 624)) + (wbMult(629) & wbMult(629 downto 627));
      v.Lvl1(423 downto 420) := (wbMult(632) & wbMult(632 downto 630)) + (wbMult(635) & wbMult(635 downto 633));
      v.Lvl1(427 downto 424) := (wbMult(638) & wbMult(638 downto 636)) + (wbMult(641) & wbMult(641 downto 639));
      v.Lvl1(431 downto 428) := (wbMult(644) & wbMult(644 downto 642)) + (wbMult(647) & wbMult(647 downto 645));
      v.Lvl1(435 downto 432) := (wbMult(650) & wbMult(650 downto 648)) + (wbMult(653) & wbMult(653 downto 651));
      v.Lvl1(439 downto 436) := (wbMult(656) & wbMult(656 downto 654)) + (wbMult(659) & wbMult(659 downto 657));
      v.Lvl1(443 downto 440) := (wbMult(662) & wbMult(662 downto 660)) + (wbMult(665) & wbMult(665 downto 663));
      v.Lvl1(447 downto 444) := (wbMult(668) & wbMult(668 downto 666)) + (wbMult(671) & wbMult(671 downto 669));
      v.Lvl1(451 downto 448) := (wbMult(674) & wbMult(674 downto 672)) + (wbMult(677) & wbMult(677 downto 675));
      v.Lvl1(455 downto 452) := (wbMult(680) & wbMult(680 downto 678)) + (wbMult(683) & wbMult(683 downto 681));
      v.Lvl1(459 downto 456) := (wbMult(686) & wbMult(686 downto 684)) + (wbMult(689) & wbMult(689 downto 687));
      v.Lvl1(463 downto 460) := (wbMult(692) & wbMult(692 downto 690)) + (wbMult(695) & wbMult(695 downto 693));
      v.Lvl1(467 downto 464) := (wbMult(698) & wbMult(698 downto 696)) + (wbMult(701) & wbMult(701 downto 699));
      v.Lvl1(471 downto 468) := (wbMult(704) & wbMult(704 downto 702)) + (wbMult(707) & wbMult(707 downto 705));
      v.Lvl1(475 downto 472) := (wbMult(710) & wbMult(710 downto 708)) + (wbMult(713) & wbMult(713 downto 711));
      v.Lvl1(479 downto 476) := (wbMult(716) & wbMult(716 downto 714)) + (wbMult(719) & wbMult(719 downto 717));
      v.Lvl1(483 downto 480) := (wbMult(722) & wbMult(722 downto 720)) + (wbMult(725) & wbMult(725 downto 723));
      v.Lvl1(487 downto 484) := (wbMult(728) & wbMult(728 downto 726)) + (wbMult(731) & wbMult(731 downto 729));
      v.Lvl1(491 downto 488) := (wbMult(734) & wbMult(734 downto 732)) + (wbMult(737) & wbMult(737 downto 735));
      v.Lvl1(495 downto 492) := (wbMult(740) & wbMult(740 downto 738)) + (wbMult(743) & wbMult(743 downto 741));
      v.Lvl1(499 downto 496) := (wbMult(746) & wbMult(746 downto 744)) + (wbMult(749) & wbMult(749 downto 747));
      v.Lvl1(503 downto 500) := (wbMult(752) & wbMult(752 downto 750)) + (wbMult(755) & wbMult(755 downto 753));
      v.Lvl1(507 downto 504) := (wbMult(758) & wbMult(758 downto 756)) + (wbMult(761) & wbMult(761 downto 759));
      v.Lvl1(511 downto 508) := (wbMult(764) & wbMult(764 downto 762)) + (wbMult(767) & wbMult(767 downto 765));
      v.Lvl1(515 downto 512) := (wbMult(770) & wbMult(770 downto 768)) + (wbMult(773) & wbMult(773 downto 771));
      v.Lvl1(519 downto 516) := (wbMult(776) & wbMult(776 downto 774)) + (wbMult(779) & wbMult(779 downto 777));
      v.Lvl1(523 downto 520) := (wbMult(782) & wbMult(782 downto 780)) + (wbMult(785) & wbMult(785 downto 783));
      v.Lvl1(527 downto 524) := (wbMult(788) & wbMult(788 downto 786)) + (wbMult(791) & wbMult(791 downto 789));
      v.Lvl1(531 downto 528) := (wbMult(794) & wbMult(794 downto 792)) + (wbMult(797) & wbMult(797 downto 795));
      v.Lvl1(535 downto 532) := (wbMult(800) & wbMult(800 downto 798)) + (wbMult(803) & wbMult(803 downto 801));
      v.Lvl1(539 downto 536) := (wbMult(806) & wbMult(806 downto 804)) + (wbMult(809) & wbMult(809 downto 807));
      v.Lvl1(543 downto 540) := (wbMult(812) & wbMult(812 downto 810)) + (wbMult(815) & wbMult(815 downto 813));
      v.Lvl1(547 downto 544) := (wbMult(818) & wbMult(818 downto 816)) + (wbMult(821) & wbMult(821 downto 819));
      v.Lvl1(551 downto 548) := (wbMult(824) & wbMult(824 downto 822)) + (wbMult(827) & wbMult(827 downto 825));
      v.Lvl1(555 downto 552) := (wbMult(830) & wbMult(830 downto 828)) + (wbMult(833) & wbMult(833 downto 831));
      v.Lvl1(559 downto 556) := (wbMult(836) & wbMult(836 downto 834)) + (wbMult(839) & wbMult(839 downto 837));
      v.Lvl1(563 downto 560) := (wbMult(842) & wbMult(842 downto 840)) + (wbMult(845) & wbMult(845 downto 843));
      v.Lvl1(567 downto 564) := (wbMult(848) & wbMult(848 downto 846)) + (wbMult(851) & wbMult(851 downto 849));
      v.Lvl1(571 downto 568) := (wbMult(854) & wbMult(854 downto 852)) + (wbMult(857) & wbMult(857 downto 855));
      v.Lvl1(575 downto 572) := (wbMult(860) & wbMult(860 downto 858)) + (wbMult(863) & wbMult(863 downto 861));
      v.Lvl1(579 downto 576) := (wbMult(866) & wbMult(866 downto 864)) + (wbMult(869) & wbMult(869 downto 867));
      v.Lvl1(583 downto 580) := (wbMult(872) & wbMult(872 downto 870)) + (wbMult(875) & wbMult(875 downto 873));
      v.Lvl1(587 downto 584) := (wbMult(878) & wbMult(878 downto 876)) + (wbMult(881) & wbMult(881 downto 879));
      v.Lvl1(591 downto 588) := (wbMult(884) & wbMult(884 downto 882)) + (wbMult(887) & wbMult(887 downto 885));
      v.Lvl1(595 downto 592) := (wbMult(890) & wbMult(890 downto 888)) + (wbMult(893) & wbMult(893 downto 891));
      v.Lvl1(599 downto 596) := (wbMult(896) & wbMult(896 downto 894)) + (wbMult(899) & wbMult(899 downto 897));
      v.Lvl1(603 downto 600) := (wbMult(902) & wbMult(902 downto 900)) + (wbMult(905) & wbMult(905 downto 903));
      v.Lvl1(607 downto 604) := (wbMult(908) & wbMult(908 downto 906)) + (wbMult(911) & wbMult(911 downto 909));
      v.Lvl1(611 downto 608) := (wbMult(914) & wbMult(914 downto 912)) + (wbMult(917) & wbMult(917 downto 915));
      v.Lvl1(615 downto 612) := (wbMult(920) & wbMult(920 downto 918)) + (wbMult(923) & wbMult(923 downto 921));
      v.Lvl1(619 downto 616) := (wbMult(926) & wbMult(926 downto 924)) + (wbMult(929) & wbMult(929 downto 927));
      v.Lvl1(623 downto 620) := (wbMult(932) & wbMult(932 downto 930)) + (wbMult(935) & wbMult(935 downto 933));
      v.Lvl1(627 downto 624) := (wbMult(938) & wbMult(938 downto 936)) + (wbMult(941) & wbMult(941 downto 939));
      v.Lvl1(631 downto 628) := (wbMult(944) & wbMult(944 downto 942)) + (wbMult(947) & wbMult(947 downto 945));
      v.Lvl1(635 downto 632) := (wbMult(950) & wbMult(950 downto 948)) + (wbMult(953) & wbMult(953 downto 951));
      v.Lvl1(639 downto 636) := (wbMult(956) & wbMult(956 downto 954)) + (wbMult(959) & wbMult(959 downto 957));
      v.Lvl1(643 downto 640) := (wbMult(962) & wbMult(962 downto 960)) + (wbMult(965) & wbMult(965 downto 963));
      v.Lvl1(647 downto 644) := (wbMult(968) & wbMult(968 downto 966)) + (wbMult(971) & wbMult(971 downto 969));
      v.Lvl1(651 downto 648) := (wbMult(974) & wbMult(974 downto 972)) + (wbMult(977) & wbMult(977 downto 975));
      v.Lvl1(655 downto 652) := (wbMult(980) & wbMult(980 downto 978)) + (wbMult(983) & wbMult(983 downto 981));
      v.Lvl1(659 downto 656) := (wbMult(986) & wbMult(986 downto 984)) + (wbMult(989) & wbMult(989 downto 987));
      v.Lvl1(663 downto 660) := (wbMult(992) & wbMult(992 downto 990)) + (wbMult(995) & wbMult(995 downto 993));
      v.Lvl1(667 downto 664) := (wbMult(998) & wbMult(998 downto 996)) + (wbMult(1001) & wbMult(1001 downto 999));
      v.Lvl1(671 downto 668) := (wbMult(1004) & wbMult(1004 downto 1002)) + (wbMult(1007) & wbMult(1007 downto 1005));
      v.Lvl1(675 downto 672) := (wbMult(1010) & wbMult(1010 downto 1008)) + (wbMult(1013) & wbMult(1013 downto 1011));
      v.Lvl1(679 downto 676) := (wbMult(1016) & wbMult(1016 downto 1014)) + (wbMult(1019) & wbMult(1019 downto 1017));
      v.Lvl1(683 downto 680) := (wbMult(1022) & wbMult(1022 downto 1020)) + (wbMult(1025) & wbMult(1025 downto 1023));
      v.Lvl1(687 downto 684) := (wbMult(1028) & wbMult(1028 downto 1026)) + (wbMult(1031) & wbMult(1031 downto 1029));
      v.Lvl1(691 downto 688) := (wbMult(1034) & wbMult(1034 downto 1032)) + (wbMult(1037) & wbMult(1037 downto 1035));
      v.Lvl1(695 downto 692) := (wbMult(1040) & wbMult(1040 downto 1038)) + (wbMult(1043) & wbMult(1043 downto 1041));
      v.Lvl1(699 downto 696) := (wbMult(1046) & wbMult(1046 downto 1044)) + (wbMult(1049) & wbMult(1049 downto 1047));
      v.Lvl1(703 downto 700) := (wbMult(1052) & wbMult(1052 downto 1050)) + (wbMult(1055) & wbMult(1055 downto 1053));
      v.Lvl1(707 downto 704) := (wbMult(1058) & wbMult(1058 downto 1056)) + (wbMult(1061) & wbMult(1061 downto 1059));
      v.Lvl1(711 downto 708) := (wbMult(1064) & wbMult(1064 downto 1062)) + (wbMult(1067) & wbMult(1067 downto 1065));
      v.Lvl1(715 downto 712) := (wbMult(1070) & wbMult(1070 downto 1068)) + (wbMult(1073) & wbMult(1073 downto 1071));
      v.Lvl1(719 downto 716) := (wbMult(1076) & wbMult(1076 downto 1074)) + (wbMult(1079) & wbMult(1079 downto 1077));
      v.Lvl1(723 downto 720) := (wbMult(1082) & wbMult(1082 downto 1080)) + (wbMult(1085) & wbMult(1085 downto 1083));
      v.Lvl1(727 downto 724) := (wbMult(1088) & wbMult(1088 downto 1086)) + (wbMult(1091) & wbMult(1091 downto 1089));
      v.Lvl1(731 downto 728) := (wbMult(1094) & wbMult(1094 downto 1092)) + (wbMult(1097) & wbMult(1097 downto 1095));
      v.Lvl1(735 downto 732) := (wbMult(1100) & wbMult(1100 downto 1098)) + (wbMult(1103) & wbMult(1103 downto 1101));
      v.Lvl1(739 downto 736) := (wbMult(1106) & wbMult(1106 downto 1104)) + (wbMult(1109) & wbMult(1109 downto 1107));
      v.Lvl1(743 downto 740) := (wbMult(1112) & wbMult(1112 downto 1110)) + (wbMult(1115) & wbMult(1115 downto 1113));
      v.Lvl1(747 downto 744) := (wbMult(1118) & wbMult(1118 downto 1116)) + (wbMult(1121) & wbMult(1121 downto 1119));
      v.Lvl1(751 downto 748) := (wbMult(1124) & wbMult(1124 downto 1122)) + (wbMult(1127) & wbMult(1127 downto 1125));
      v.Lvl1(755 downto 752) := (wbMult(1130) & wbMult(1130 downto 1128)) + (wbMult(1133) & wbMult(1133 downto 1131));
      v.Lvl1(759 downto 756) := (wbMult(1136) & wbMult(1136 downto 1134)) + (wbMult(1139) & wbMult(1139 downto 1137));
      v.Lvl1(763 downto 760) := (wbMult(1142) & wbMult(1142 downto 1140)) + (wbMult(1145) & wbMult(1145 downto 1143));
      v.Lvl1(767 downto 764) := (wbMult(1148) & wbMult(1148 downto 1146)) + (wbMult(1151) & wbMult(1151 downto 1149));
      v.Lvl1(771 downto 768) := (wbMult(1154) & wbMult(1154 downto 1152)) + (wbMult(1157) & wbMult(1157 downto 1155));
      v.Lvl1(775 downto 772) := (wbMult(1160) & wbMult(1160 downto 1158)) + (wbMult(1163) & wbMult(1163 downto 1161));
      v.Lvl1(779 downto 776) := (wbMult(1166) & wbMult(1166 downto 1164)) + (wbMult(1169) & wbMult(1169 downto 1167));
      v.Lvl1(783 downto 780) := (wbMult(1172) & wbMult(1172 downto 1170)) + (wbMult(1175) & wbMult(1175 downto 1173));
      v.Lvl1(787 downto 784) := (wbMult(1178) & wbMult(1178 downto 1176)) + (wbMult(1181) & wbMult(1181 downto 1179));
      v.Lvl1(791 downto 788) := (wbMult(1184) & wbMult(1184 downto 1182)) + (wbMult(1187) & wbMult(1187 downto 1185));
      v.Lvl1(795 downto 792) := (wbMult(1190) & wbMult(1190 downto 1188)) + (wbMult(1193) & wbMult(1193 downto 1191));
      v.Lvl1(799 downto 796) := (wbMult(1196) & wbMult(1196 downto 1194)) + (wbMult(1199) & wbMult(1199 downto 1197));
      v.Lvl1(803 downto 800) := (wbMult(1202) & wbMult(1202 downto 1200)) + (wbMult(1205) & wbMult(1205 downto 1203));
      v.Lvl1(807 downto 804) := (wbMult(1208) & wbMult(1208 downto 1206)) + (wbMult(1211) & wbMult(1211 downto 1209));
      v.Lvl1(811 downto 808) := (wbMult(1214) & wbMult(1214 downto 1212)) + (wbMult(1217) & wbMult(1217 downto 1215));
      v.Lvl1(815 downto 812) := (wbMult(1220) & wbMult(1220 downto 1218)) + (wbMult(1223) & wbMult(1223 downto 1221));
      v.Lvl1(819 downto 816) := (wbMult(1226) & wbMult(1226 downto 1224)) + (wbMult(1229) & wbMult(1229 downto 1227));
      v.Lvl1(823 downto 820) := (wbMult(1232) & wbMult(1232 downto 1230)) + (wbMult(1235) & wbMult(1235 downto 1233));
      v.Lvl1(827 downto 824) := (wbMult(1238) & wbMult(1238 downto 1236)) + (wbMult(1241) & wbMult(1241 downto 1239));
      v.Lvl1(831 downto 828) := (wbMult(1244) & wbMult(1244 downto 1242)) + (wbMult(1247) & wbMult(1247 downto 1245));
      v.Lvl1(835 downto 832) := (wbMult(1250) & wbMult(1250 downto 1248)) + (wbMult(1253) & wbMult(1253 downto 1251));
      v.Lvl1(839 downto 836) := (wbMult(1256) & wbMult(1256 downto 1254)) + (wbMult(1259) & wbMult(1259 downto 1257));
      v.Lvl1(843 downto 840) := (wbMult(1262) & wbMult(1262 downto 1260)) + (wbMult(1265) & wbMult(1265 downto 1263));
      v.Lvl1(847 downto 844) := (wbMult(1268) & wbMult(1268 downto 1266)) + (wbMult(1271) & wbMult(1271 downto 1269));
      v.Lvl1(851 downto 848) := (wbMult(1274) & wbMult(1274 downto 1272)) + (wbMult(1277) & wbMult(1277 downto 1275));
      v.Lvl1(855 downto 852) := (wbMult(1280) & wbMult(1280 downto 1278)) + (wbMult(1283) & wbMult(1283 downto 1281));
      v.Lvl1(859 downto 856) := (wbMult(1286) & wbMult(1286 downto 1284)) + (wbMult(1289) & wbMult(1289 downto 1287));
      v.Lvl1(863 downto 860) := (wbMult(1292) & wbMult(1292 downto 1290)) + (wbMult(1295) & wbMult(1295 downto 1293));
      v.Lvl1(867 downto 864) := (wbMult(1298) & wbMult(1298 downto 1296)) + (wbMult(1301) & wbMult(1301 downto 1299));
      v.Lvl1(871 downto 868) := (wbMult(1304) & wbMult(1304 downto 1302)) + (wbMult(1307) & wbMult(1307 downto 1305));
      v.Lvl1(875 downto 872) := (wbMult(1310) & wbMult(1310 downto 1308)) + (wbMult(1313) & wbMult(1313 downto 1311));
      v.Lvl1(879 downto 876) := (wbMult(1316) & wbMult(1316 downto 1314)) + (wbMult(1319) & wbMult(1319 downto 1317));
      v.Lvl1(883 downto 880) := (wbMult(1322) & wbMult(1322 downto 1320)) + (wbMult(1325) & wbMult(1325 downto 1323));
      v.Lvl1(887 downto 884) := (wbMult(1328) & wbMult(1328 downto 1326)) + (wbMult(1331) & wbMult(1331 downto 1329));
      v.Lvl1(891 downto 888) := (wbMult(1334) & wbMult(1334 downto 1332)) + (wbMult(1337) & wbMult(1337 downto 1335));
      v.Lvl1(895 downto 892) := (wbMult(1340) & wbMult(1340 downto 1338)) + (wbMult(1343) & wbMult(1343 downto 1341));
      v.Lvl1(899 downto 896) := (wbMult(1346) & wbMult(1346 downto 1344)) + (wbMult(1349) & wbMult(1349 downto 1347));
      v.Lvl1(903 downto 900) := (wbMult(1352) & wbMult(1352 downto 1350)) + (wbMult(1355) & wbMult(1355 downto 1353));
      v.Lvl1(907 downto 904) := (wbMult(1358) & wbMult(1358 downto 1356)) + (wbMult(1361) & wbMult(1361 downto 1359));
      v.Lvl1(911 downto 908) := (wbMult(1364) & wbMult(1364 downto 1362)) + (wbMult(1367) & wbMult(1367 downto 1365));
      v.Lvl1(915 downto 912) := (wbMult(1370) & wbMult(1370 downto 1368)) + (wbMult(1373) & wbMult(1373 downto 1371));
      v.Lvl1(919 downto 916) := (wbMult(1376) & wbMult(1376 downto 1374)) + (wbMult(1379) & wbMult(1379 downto 1377));
      v.Lvl1(923 downto 920) := (wbMult(1382) & wbMult(1382 downto 1380)) + (wbMult(1385) & wbMult(1385 downto 1383));
      v.Lvl1(927 downto 924) := (wbMult(1388) & wbMult(1388 downto 1386)) + (wbMult(1391) & wbMult(1391 downto 1389));
      v.Lvl1(931 downto 928) := (wbMult(1394) & wbMult(1394 downto 1392)) + (wbMult(1397) & wbMult(1397 downto 1395));
      v.Lvl1(935 downto 932) := (wbMult(1400) & wbMult(1400 downto 1398)) + (wbMult(1403) & wbMult(1403 downto 1401));
      v.Lvl1(939 downto 936) := (wbMult(1406) & wbMult(1406 downto 1404)) + (wbMult(1409) & wbMult(1409 downto 1407));
      v.Lvl1(943 downto 940) := (wbMult(1412) & wbMult(1412 downto 1410)) + (wbMult(1415) & wbMult(1415 downto 1413));
      v.Lvl1(947 downto 944) := (wbMult(1418) & wbMult(1418 downto 1416)) + (wbMult(1421) & wbMult(1421 downto 1419));
      v.Lvl1(951 downto 948) := (wbMult(1424) & wbMult(1424 downto 1422)) + (wbMult(1427) & wbMult(1427 downto 1425));
      v.Lvl1(955 downto 952) := (wbMult(1430) & wbMult(1430 downto 1428)) + (wbMult(1433) & wbMult(1433 downto 1431));
      v.Lvl1(959 downto 956) := (wbMult(1436) & wbMult(1436 downto 1434)) + (wbMult(1439) & wbMult(1439 downto 1437));
      v.Lvl1(963 downto 960) := (wbMult(1442) & wbMult(1442 downto 1440)) + (wbMult(1445) & wbMult(1445 downto 1443));
      v.Lvl1(967 downto 964) := (wbMult(1448) & wbMult(1448 downto 1446)) + (wbMult(1451) & wbMult(1451 downto 1449));
      v.Lvl1(971 downto 968) := (wbMult(1454) & wbMult(1454 downto 1452)) + (wbMult(1457) & wbMult(1457 downto 1455));
      v.Lvl1(975 downto 972) := (wbMult(1460) & wbMult(1460 downto 1458)) + (wbMult(1463) & wbMult(1463 downto 1461));
      v.Lvl1(979 downto 976) := (wbMult(1466) & wbMult(1466 downto 1464)) + (wbMult(1469) & wbMult(1469 downto 1467));
      v.Lvl1(983 downto 980) := (wbMult(1472) & wbMult(1472 downto 1470)) + (wbMult(1475) & wbMult(1475 downto 1473));
      v.Lvl1(987 downto 984) := (wbMult(1478) & wbMult(1478 downto 1476)) + (wbMult(1481) & wbMult(1481 downto 1479));
      v.Lvl1(991 downto 988) := (wbMult(1484) & wbMult(1484 downto 1482)) + (wbMult(1487) & wbMult(1487 downto 1485));
      v.Lvl1(995 downto 992) := (wbMult(1490) & wbMult(1490 downto 1488)) + (wbMult(1493) & wbMult(1493 downto 1491));
      v.Lvl1(999 downto 996) := (wbMult(1496) & wbMult(1496 downto 1494)) + (wbMult(1499) & wbMult(1499 downto 1497));
      v.Lvl1(1003 downto 1000) := (wbMult(1502) & wbMult(1502 downto 1500)) + (wbMult(1505) & wbMult(1505 downto 1503));
      v.Lvl1(1007 downto 1004) := (wbMult(1508) & wbMult(1508 downto 1506)) + (wbMult(1511) & wbMult(1511 downto 1509));
      v.Lvl1(1011 downto 1008) := (wbMult(1514) & wbMult(1514 downto 1512)) + (wbMult(1517) & wbMult(1517 downto 1515));
      v.Lvl1(1015 downto 1012) := (wbMult(1520) & wbMult(1520 downto 1518)) + (wbMult(1523) & wbMult(1523 downto 1521));
      v.Lvl1(1019 downto 1016) := (wbMult(1526) & wbMult(1526 downto 1524)) + (wbMult(1529) & wbMult(1529 downto 1527));
      v.Lvl1(1023 downto 1020) := (wbMult(1532) & wbMult(1532 downto 1530)) + (wbMult(1535) & wbMult(1535 downto 1533));
      v.Lvl1(1027 downto 1024) := (wbMult(1538) & wbMult(1538 downto 1536)) + (wbMult(1541) & wbMult(1541 downto 1539));
      v.Lvl1(1031 downto 1028) := (wbMult(1544) & wbMult(1544 downto 1542)) + (wbMult(1547) & wbMult(1547 downto 1545));
      v.Lvl1(1035 downto 1032) := (wbMult(1550) & wbMult(1550 downto 1548)) + (wbMult(1553) & wbMult(1553 downto 1551));
      v.Lvl1(1039 downto 1036) := (wbMult(1556) & wbMult(1556 downto 1554)) + (wbMult(1559) & wbMult(1559 downto 1557));
      v.Lvl1(1043 downto 1040) := (wbMult(1562) & wbMult(1562 downto 1560)) + (wbMult(1565) & wbMult(1565 downto 1563));
      v.Lvl1(1047 downto 1044) := (wbMult(1568) & wbMult(1568 downto 1566)) + (wbMult(1571) & wbMult(1571 downto 1569));
      v.Lvl1(1051 downto 1048) := (wbMult(1574) & wbMult(1574 downto 1572)) + (wbMult(1577) & wbMult(1577 downto 1575));
      v.Lvl1(1055 downto 1052) := (wbMult(1580) & wbMult(1580 downto 1578)) + (wbMult(1583) & wbMult(1583 downto 1581));
      v.Lvl1(1059 downto 1056) := (wbMult(1586) & wbMult(1586 downto 1584)) + (wbMult(1589) & wbMult(1589 downto 1587));
      v.Lvl1(1063 downto 1060) := (wbMult(1592) & wbMult(1592 downto 1590)) + (wbMult(1595) & wbMult(1595 downto 1593));
      v.Lvl1(1067 downto 1064) := (wbMult(1598) & wbMult(1598 downto 1596)) + (wbMult(1601) & wbMult(1601 downto 1599));
      v.Lvl1(1071 downto 1068) := (wbMult(1604) & wbMult(1604 downto 1602)) + (wbMult(1607) & wbMult(1607 downto 1605));
      v.Lvl1(1075 downto 1072) := (wbMult(1610) & wbMult(1610 downto 1608)) + (wbMult(1613) & wbMult(1613 downto 1611));
      v.Lvl1(1079 downto 1076) := (wbMult(1616) & wbMult(1616 downto 1614)) + (wbMult(1619) & wbMult(1619 downto 1617));
      v.Lvl1(1083 downto 1080) := (wbMult(1622) & wbMult(1622 downto 1620)) + (wbMult(1625) & wbMult(1625 downto 1623));
      v.Lvl1(1087 downto 1084) := (wbMult(1628) & wbMult(1628 downto 1626)) + (wbMult(1631) & wbMult(1631 downto 1629));
      v.Lvl1(1091 downto 1088) := (wbMult(1634) & wbMult(1634 downto 1632)) + (wbMult(1637) & wbMult(1637 downto 1635));
      v.Lvl1(1095 downto 1092) := (wbMult(1640) & wbMult(1640 downto 1638)) + (wbMult(1643) & wbMult(1643 downto 1641));
      v.Lvl1(1099 downto 1096) := (wbMult(1646) & wbMult(1646 downto 1644)) + (wbMult(1649) & wbMult(1649 downto 1647));
      v.Lvl1(1103 downto 1100) := (wbMult(1652) & wbMult(1652 downto 1650)) + (wbMult(1655) & wbMult(1655 downto 1653));
      v.Lvl1(1107 downto 1104) := (wbMult(1658) & wbMult(1658 downto 1656)) + (wbMult(1661) & wbMult(1661 downto 1659));
      v.Lvl1(1111 downto 1108) := (wbMult(1664) & wbMult(1664 downto 1662)) + (wbMult(1667) & wbMult(1667 downto 1665));
      v.Lvl1(1115 downto 1112) := (wbMult(1670) & wbMult(1670 downto 1668)) + (wbMult(1673) & wbMult(1673 downto 1671));
      v.Lvl1(1119 downto 1116) := (wbMult(1676) & wbMult(1676 downto 1674)) + (wbMult(1679) & wbMult(1679 downto 1677));
      v.Lvl1(1123 downto 1120) := (wbMult(1682) & wbMult(1682 downto 1680)) + (wbMult(1685) & wbMult(1685 downto 1683));
      v.Lvl1(1127 downto 1124) := (wbMult(1688) & wbMult(1688 downto 1686)) + (wbMult(1691) & wbMult(1691 downto 1689));
      v.Lvl1(1131 downto 1128) := (wbMult(1694) & wbMult(1694 downto 1692)) + (wbMult(1697) & wbMult(1697 downto 1695));
      v.Lvl1(1135 downto 1132) := (wbMult(1700) & wbMult(1700 downto 1698)) + (wbMult(1703) & wbMult(1703 downto 1701));
      v.Lvl1(1139 downto 1136) := (wbMult(1706) & wbMult(1706 downto 1704)) + (wbMult(1709) & wbMult(1709 downto 1707));
      v.Lvl1(1143 downto 1140) := (wbMult(1712) & wbMult(1712 downto 1710)) + (wbMult(1715) & wbMult(1715 downto 1713));
      v.Lvl1(1147 downto 1144) := (wbMult(1718) & wbMult(1718 downto 1716)) + (wbMult(1721) & wbMult(1721 downto 1719));
      v.Lvl1(1151 downto 1148) := (wbMult(1724) & wbMult(1724 downto 1722)) + (wbMult(1727) & wbMult(1727 downto 1725));
      v.Lvl1(1155 downto 1152) := (wbMult(1730) & wbMult(1730 downto 1728)) + (wbMult(1733) & wbMult(1733 downto 1731));
      v.Lvl1(1159 downto 1156) := (wbMult(1736) & wbMult(1736 downto 1734)) + (wbMult(1739) & wbMult(1739 downto 1737));
      v.Lvl1(1163 downto 1160) := (wbMult(1742) & wbMult(1742 downto 1740)) + (wbMult(1745) & wbMult(1745 downto 1743));
      v.Lvl1(1167 downto 1164) := (wbMult(1748) & wbMult(1748 downto 1746)) + (wbMult(1751) & wbMult(1751 downto 1749));
      v.Lvl1(1171 downto 1168) := (wbMult(1754) & wbMult(1754 downto 1752)) + (wbMult(1757) & wbMult(1757 downto 1755));
      v.Lvl1(1175 downto 1172) := (wbMult(1760) & wbMult(1760 downto 1758)) + (wbMult(1763) & wbMult(1763 downto 1761));
      v.Lvl1(1179 downto 1176) := (wbMult(1766) & wbMult(1766 downto 1764)) + (wbMult(1769) & wbMult(1769 downto 1767));
      v.Lvl1(1183 downto 1180) := (wbMult(1772) & wbMult(1772 downto 1770)) + (wbMult(1775) & wbMult(1775 downto 1773));
      v.Lvl1(1187 downto 1184) := (wbMult(1778) & wbMult(1778 downto 1776)) + (wbMult(1781) & wbMult(1781 downto 1779));
      v.Lvl1(1191 downto 1188) := (wbMult(1784) & wbMult(1784 downto 1782)) + (wbMult(1787) & wbMult(1787 downto 1785));
      v.Lvl1(1195 downto 1192) := (wbMult(1790) & wbMult(1790 downto 1788)) + (wbMult(1793) & wbMult(1793 downto 1791));
      v.Lvl1(1199 downto 1196) := (wbMult(1796) & wbMult(1796 downto 1794)) + (wbMult(1799) & wbMult(1799 downto 1797));
      v.Lvl1(1203 downto 1200) := (wbMult(1802) & wbMult(1802 downto 1800)) + (wbMult(1805) & wbMult(1805 downto 1803));
      v.Lvl1(1207 downto 1204) := (wbMult(1808) & wbMult(1808 downto 1806)) + (wbMult(1811) & wbMult(1811 downto 1809));
      v.Lvl1(1211 downto 1208) := (wbMult(1814) & wbMult(1814 downto 1812)) + (wbMult(1817) & wbMult(1817 downto 1815));
      v.Lvl1(1215 downto 1212) := (wbMult(1820) & wbMult(1820 downto 1818)) + (wbMult(1823) & wbMult(1823 downto 1821));
      v.Lvl1(1219 downto 1216) := (wbMult(1826) & wbMult(1826 downto 1824)) + (wbMult(1829) & wbMult(1829 downto 1827));
      v.Lvl1(1223 downto 1220) := (wbMult(1832) & wbMult(1832 downto 1830)) + (wbMult(1835) & wbMult(1835 downto 1833));
      v.Lvl1(1227 downto 1224) := (wbMult(1838) & wbMult(1838 downto 1836)) + (wbMult(1841) & wbMult(1841 downto 1839));
      v.Lvl1(1231 downto 1228) := (wbMult(1844) & wbMult(1844 downto 1842)) + (wbMult(1847) & wbMult(1847 downto 1845));
      v.Lvl1(1235 downto 1232) := (wbMult(1850) & wbMult(1850 downto 1848)) + (wbMult(1853) & wbMult(1853 downto 1851));
      v.Lvl1(1239 downto 1236) := (wbMult(1856) & wbMult(1856 downto 1854)) + (wbMult(1859) & wbMult(1859 downto 1857));
      v.Lvl1(1243 downto 1240) := (wbMult(1862) & wbMult(1862 downto 1860)) + (wbMult(1865) & wbMult(1865 downto 1863));
      v.Lvl1(1247 downto 1244) := (wbMult(1868) & wbMult(1868 downto 1866)) + (wbMult(1871) & wbMult(1871 downto 1869));
      v.Lvl1(1251 downto 1248) := (wbMult(1874) & wbMult(1874 downto 1872)) + (wbMult(1877) & wbMult(1877 downto 1875));
      v.Lvl1(1255 downto 1252) := (wbMult(1880) & wbMult(1880 downto 1878)) + (wbMult(1883) & wbMult(1883 downto 1881));
      v.Lvl1(1259 downto 1256) := (wbMult(1886) & wbMult(1886 downto 1884)) + (wbMult(1889) & wbMult(1889 downto 1887));
      v.Lvl1(1263 downto 1260) := (wbMult(1892) & wbMult(1892 downto 1890)) + (wbMult(1895) & wbMult(1895 downto 1893));
      v.Lvl1(1267 downto 1264) := (wbMult(1898) & wbMult(1898 downto 1896)) + (wbMult(1901) & wbMult(1901 downto 1899));
      v.Lvl1(1271 downto 1268) := (wbMult(1904) & wbMult(1904 downto 1902)) + (wbMult(1907) & wbMult(1907 downto 1905));
      v.Lvl1(1275 downto 1272) := (wbMult(1910) & wbMult(1910 downto 1908)) + (wbMult(1913) & wbMult(1913 downto 1911));
      v.Lvl1(1279 downto 1276) := (wbMult(1916) & wbMult(1916 downto 1914)) + (wbMult(1919) & wbMult(1919 downto 1917));
      v.Lvl1(1283 downto 1280) := (wbMult(1922) & wbMult(1922 downto 1920)) + (wbMult(1925) & wbMult(1925 downto 1923));
      v.Lvl1(1287 downto 1284) := (wbMult(1928) & wbMult(1928 downto 1926)) + (wbMult(1931) & wbMult(1931 downto 1929));
      v.Lvl1(1291 downto 1288) := (wbMult(1934) & wbMult(1934 downto 1932)) + (wbMult(1937) & wbMult(1937 downto 1935));
      v.Lvl1(1295 downto 1292) := (wbMult(1940) & wbMult(1940 downto 1938)) + (wbMult(1943) & wbMult(1943 downto 1941));
      v.Lvl1(1299 downto 1296) := (wbMult(1946) & wbMult(1946 downto 1944)) + (wbMult(1949) & wbMult(1949 downto 1947));
      v.Lvl1(1303 downto 1300) := (wbMult(1952) & wbMult(1952 downto 1950)) + (wbMult(1955) & wbMult(1955 downto 1953));
      v.Lvl1(1307 downto 1304) := (wbMult(1958) & wbMult(1958 downto 1956)) + (wbMult(1961) & wbMult(1961 downto 1959));
      v.Lvl1(1311 downto 1308) := (wbMult(1964) & wbMult(1964 downto 1962)) + (wbMult(1967) & wbMult(1967 downto 1965));
      v.Lvl1(1315 downto 1312) := (wbMult(1970) & wbMult(1970 downto 1968)) + (wbMult(1973) & wbMult(1973 downto 1971));
      v.Lvl1(1319 downto 1316) := (wbMult(1976) & wbMult(1976 downto 1974)) + (wbMult(1979) & wbMult(1979 downto 1977));
      v.Lvl1(1323 downto 1320) := (wbMult(1982) & wbMult(1982 downto 1980)) + (wbMult(1985) & wbMult(1985 downto 1983));
      v.Lvl1(1327 downto 1324) := (wbMult(1988) & wbMult(1988 downto 1986)) + (wbMult(1991) & wbMult(1991 downto 1989));
      v.Lvl1(1331 downto 1328) := (wbMult(1994) & wbMult(1994 downto 1992)) + (wbMult(1997) & wbMult(1997 downto 1995));
      v.Lvl1(1335 downto 1332) := (wbMult(2000) & wbMult(2000 downto 1998)) + (wbMult(2003) & wbMult(2003 downto 2001));
      v.Lvl1(1339 downto 1336) := (wbMult(2006) & wbMult(2006 downto 2004)) + (wbMult(2009) & wbMult(2009 downto 2007));
      v.Lvl1(1343 downto 1340) := (wbMult(2012) & wbMult(2012 downto 2010)) + (wbMult(2015) & wbMult(2015 downto 2013));
      v.Lvl1(1347 downto 1344) := (wbMult(2018) & wbMult(2018 downto 2016)) + (wbMult(2021) & wbMult(2021 downto 2019));
      v.Lvl1(1351 downto 1348) := (wbMult(2024) & wbMult(2024 downto 2022)) + (wbMult(2027) & wbMult(2027 downto 2025));
      v.Lvl1(1355 downto 1352) := (wbMult(2030) & wbMult(2030 downto 2028)) + (wbMult(2033) & wbMult(2033 downto 2031));
      v.Lvl1(1359 downto 1356) := (wbMult(2036) & wbMult(2036 downto 2034)) + (wbMult(2039) & wbMult(2039 downto 2037));
      v.Lvl1(1363 downto 1360) := (wbMult(2042) & wbMult(2042 downto 2040)) + (wbMult(2045) & wbMult(2045 downto 2043));
      v.Lvl1(1367 downto 1364) := (wbMult(2048) & wbMult(2048 downto 2046)) + (wbMult(2051) & wbMult(2051 downto 2049));
      v.Lvl1(1371 downto 1368) := (wbMult(2054) & wbMult(2054 downto 2052)) + (wbMult(2057) & wbMult(2057 downto 2055));
      v.Lvl1(1375 downto 1372) := (wbMult(2060) & wbMult(2060 downto 2058)) + (wbMult(2063) & wbMult(2063 downto 2061));
      v.Lvl1(1379 downto 1376) := (wbMult(2066) & wbMult(2066 downto 2064)) + (wbMult(2069) & wbMult(2069 downto 2067));
      v.Lvl1(1383 downto 1380) := (wbMult(2072) & wbMult(2072 downto 2070)) + (wbMult(2075) & wbMult(2075 downto 2073));
      v.Lvl1(1387 downto 1384) := (wbMult(2078) & wbMult(2078 downto 2076)) + (wbMult(2081) & wbMult(2081 downto 2079));
      v.Lvl1(1391 downto 1388) := (wbMult(2084) & wbMult(2084 downto 2082)) + (wbMult(2087) & wbMult(2087 downto 2085));
      v.Lvl1(1395 downto 1392) := (wbMult(2090) & wbMult(2090 downto 2088)) + (wbMult(2093) & wbMult(2093 downto 2091));
      v.Lvl1(1399 downto 1396) := (wbMult(2096) & wbMult(2096 downto 2094)) + (wbMult(2099) & wbMult(2099 downto 2097));
      v.Lvl1(1403 downto 1400) := (wbMult(2102) & wbMult(2102 downto 2100)) + (wbMult(2105) & wbMult(2105 downto 2103));
      v.Lvl1(1407 downto 1404) := (wbMult(2108) & wbMult(2108 downto 2106)) + (wbMult(2111) & wbMult(2111 downto 2109));
      v.Lvl1(1411 downto 1408) := (wbMult(2114) & wbMult(2114 downto 2112)) + (wbMult(2117) & wbMult(2117 downto 2115));
      v.Lvl1(1415 downto 1412) := (wbMult(2120) & wbMult(2120 downto 2118)) + (wbMult(2123) & wbMult(2123 downto 2121));
      v.Lvl1(1419 downto 1416) := (wbMult(2126) & wbMult(2126 downto 2124)) + (wbMult(2129) & wbMult(2129 downto 2127));
      v.Lvl1(1423 downto 1420) := (wbMult(2132) & wbMult(2132 downto 2130)) + (wbMult(2135) & wbMult(2135 downto 2133));
      v.Lvl1(1427 downto 1424) := (wbMult(2138) & wbMult(2138 downto 2136)) + (wbMult(2141) & wbMult(2141 downto 2139));
      v.Lvl1(1431 downto 1428) := (wbMult(2144) & wbMult(2144 downto 2142)) + (wbMult(2147) & wbMult(2147 downto 2145));
      v.Lvl1(1435 downto 1432) := (wbMult(2150) & wbMult(2150 downto 2148)) + (wbMult(2153) & wbMult(2153 downto 2151));
      v.Lvl1(1439 downto 1436) := (wbMult(2156) & wbMult(2156 downto 2154)) + (wbMult(2159) & wbMult(2159 downto 2157));
      v.Lvl1(1443 downto 1440) := (wbMult(2162) & wbMult(2162 downto 2160)) + (wbMult(2165) & wbMult(2165 downto 2163));
      v.Lvl1(1447 downto 1444) := (wbMult(2168) & wbMult(2168 downto 2166)) + (wbMult(2171) & wbMult(2171 downto 2169));
      v.Lvl1(1451 downto 1448) := (wbMult(2174) & wbMult(2174 downto 2172)) + (wbMult(2177) & wbMult(2177 downto 2175));
      v.Lvl1(1455 downto 1452) := (wbMult(2180) & wbMult(2180 downto 2178)) + (wbMult(2183) & wbMult(2183 downto 2181));
      v.Lvl1(1459 downto 1456) := (wbMult(2186) & wbMult(2186 downto 2184)) + (wbMult(2189) & wbMult(2189 downto 2187));
      v.Lvl1(1463 downto 1460) := (wbMult(2192) & wbMult(2192 downto 2190)) + (wbMult(2195) & wbMult(2195 downto 2193));
      v.Lvl1(1467 downto 1464) := (wbMult(2198) & wbMult(2198 downto 2196)) + (wbMult(2201) & wbMult(2201 downto 2199));
      v.Lvl1(1471 downto 1468) := (wbMult(2204) & wbMult(2204 downto 2202)) + (wbMult(2207) & wbMult(2207 downto 2205));
      v.Lvl1(1475 downto 1472) := (wbMult(2210) & wbMult(2210 downto 2208)) + (wbMult(2213) & wbMult(2213 downto 2211));
      v.Lvl1(1479 downto 1476) := (wbMult(2216) & wbMult(2216 downto 2214)) + (wbMult(2219) & wbMult(2219 downto 2217));
      v.Lvl1(1483 downto 1480) := (wbMult(2222) & wbMult(2222 downto 2220)) + (wbMult(2225) & wbMult(2225 downto 2223));
      v.Lvl1(1487 downto 1484) := (wbMult(2228) & wbMult(2228 downto 2226)) + (wbMult(2231) & wbMult(2231 downto 2229));
      v.Lvl1(1491 downto 1488) := (wbMult(2234) & wbMult(2234 downto 2232)) + (wbMult(2237) & wbMult(2237 downto 2235));
      v.Lvl1(1495 downto 1492) := (wbMult(2240) & wbMult(2240 downto 2238)) + (wbMult(2243) & wbMult(2243 downto 2241));
      v.Lvl1(1499 downto 1496) := (wbMult(2246) & wbMult(2246 downto 2244)) + (wbMult(2249) & wbMult(2249 downto 2247));
      v.Lvl1(1503 downto 1500) := (wbMult(2252) & wbMult(2252 downto 2250)) + (wbMult(2255) & wbMult(2255 downto 2253));
      v.Lvl1(1507 downto 1504) := (wbMult(2258) & wbMult(2258 downto 2256)) + (wbMult(2261) & wbMult(2261 downto 2259));
      v.Lvl1(1511 downto 1508) := (wbMult(2264) & wbMult(2264 downto 2262)) + (wbMult(2267) & wbMult(2267 downto 2265));
      v.Lvl1(1515 downto 1512) := (wbMult(2270) & wbMult(2270 downto 2268)) + (wbMult(2273) & wbMult(2273 downto 2271));
      v.Lvl1(1519 downto 1516) := (wbMult(2276) & wbMult(2276 downto 2274)) + (wbMult(2279) & wbMult(2279 downto 2277));
      v.Lvl1(1523 downto 1520) := (wbMult(2282) & wbMult(2282 downto 2280)) + (wbMult(2285) & wbMult(2285 downto 2283));
      v.Lvl1(1527 downto 1524) := (wbMult(2288) & wbMult(2288 downto 2286)) + (wbMult(2291) & wbMult(2291 downto 2289));
      v.Lvl1(1531 downto 1528) := (wbMult(2294) & wbMult(2294 downto 2292)) + (wbMult(2297) & wbMult(2297 downto 2295));
      v.Lvl1(1535 downto 1532) := (wbMult(2300) & wbMult(2300 downto 2298)) + (wbMult(2303) & wbMult(2303 downto 2301));
      v.Lvl1(1539 downto 1536) := (wbMult(2306) & wbMult(2306 downto 2304)) + (wbMult(2309) & wbMult(2309 downto 2307));
      v.Lvl1(1543 downto 1540) := (wbMult(2312) & wbMult(2312 downto 2310)) + (wbMult(2315) & wbMult(2315 downto 2313));
      v.Lvl1(1547 downto 1544) := (wbMult(2318) & wbMult(2318 downto 2316)) + (wbMult(2321) & wbMult(2321 downto 2319));
      v.Lvl1(1551 downto 1548) := (wbMult(2324) & wbMult(2324 downto 2322)) + (wbMult(2327) & wbMult(2327 downto 2325));
      v.Lvl1(1555 downto 1552) := (wbMult(2330) & wbMult(2330 downto 2328)) + (wbMult(2333) & wbMult(2333 downto 2331));
      v.Lvl1(1559 downto 1556) := (wbMult(2336) & wbMult(2336 downto 2334)) + (wbMult(2339) & wbMult(2339 downto 2337));
      v.Lvl1(1563 downto 1560) := (wbMult(2342) & wbMult(2342 downto 2340)) + (wbMult(2345) & wbMult(2345 downto 2343));
      v.Lvl1(1567 downto 1564) := (wbMult(2348) & wbMult(2348 downto 2346)) + (wbMult(2351) & wbMult(2351 downto 2349));
      v.Lvl1(1571 downto 1568) := (wbMult(2354) & wbMult(2354 downto 2352)) + (wbMult(2357) & wbMult(2357 downto 2355));
      v.Lvl1(1575 downto 1572) := (wbMult(2360) & wbMult(2360 downto 2358)) + (wbMult(2363) & wbMult(2363 downto 2361));
      v.Lvl1(1579 downto 1576) := (wbMult(2366) & wbMult(2366 downto 2364)) + (wbMult(2369) & wbMult(2369 downto 2367));
      v.Lvl1(1583 downto 1580) := (wbMult(2372) & wbMult(2372 downto 2370)) + (wbMult(2375) & wbMult(2375 downto 2373));
      v.Lvl1(1587 downto 1584) := (wbMult(2378) & wbMult(2378 downto 2376)) + (wbMult(2381) & wbMult(2381 downto 2379));
      v.Lvl1(1591 downto 1588) := (wbMult(2384) & wbMult(2384 downto 2382)) + (wbMult(2387) & wbMult(2387 downto 2385));
      v.Lvl1(1595 downto 1592) := (wbMult(2390) & wbMult(2390 downto 2388)) + (wbMult(2393) & wbMult(2393 downto 2391));
      v.Lvl1(1599 downto 1596) := (wbMult(2396) & wbMult(2396 downto 2394)) + (wbMult(2399) & wbMult(2399 downto 2397));
      v.Lvl1(1603 downto 1600) := (wbMult(2402) & wbMult(2402 downto 2400)) + (wbMult(2405) & wbMult(2405 downto 2403));
      v.Lvl1(1607 downto 1604) := (wbMult(2408) & wbMult(2408 downto 2406)) + (wbMult(2411) & wbMult(2411 downto 2409));
      v.Lvl1(1611 downto 1608) := (wbMult(2414) & wbMult(2414 downto 2412)) + (wbMult(2417) & wbMult(2417 downto 2415));
      v.Lvl1(1615 downto 1612) := (wbMult(2420) & wbMult(2420 downto 2418)) + (wbMult(2423) & wbMult(2423 downto 2421));
      v.Lvl1(1619 downto 1616) := (wbMult(2426) & wbMult(2426 downto 2424)) + (wbMult(2429) & wbMult(2429 downto 2427));
      v.Lvl1(1623 downto 1620) := (wbMult(2432) & wbMult(2432 downto 2430)) + (wbMult(2435) & wbMult(2435 downto 2433));
      v.Lvl1(1627 downto 1624) := (wbMult(2438) & wbMult(2438 downto 2436)) + (wbMult(2441) & wbMult(2441 downto 2439));
      v.Lvl1(1631 downto 1628) := (wbMult(2444) & wbMult(2444 downto 2442)) + (wbMult(2447) & wbMult(2447 downto 2445));
      v.Lvl1(1635 downto 1632) := (wbMult(2450) & wbMult(2450 downto 2448)) + (wbMult(2453) & wbMult(2453 downto 2451));
      v.Lvl1(1639 downto 1636) := (wbMult(2456) & wbMult(2456 downto 2454)) + (wbMult(2459) & wbMult(2459 downto 2457));
      v.Lvl1(1643 downto 1640) := (wbMult(2462) & wbMult(2462 downto 2460)) + (wbMult(2465) & wbMult(2465 downto 2463));
      v.Lvl1(1647 downto 1644) := (wbMult(2468) & wbMult(2468 downto 2466)) + (wbMult(2471) & wbMult(2471 downto 2469));
      v.Lvl1(1651 downto 1648) := (wbMult(2474) & wbMult(2474 downto 2472)) + (wbMult(2477) & wbMult(2477 downto 2475));
      v.Lvl1(1655 downto 1652) := (wbMult(2480) & wbMult(2480 downto 2478)) + (wbMult(2483) & wbMult(2483 downto 2481));
      v.Lvl1(1659 downto 1656) := (wbMult(2486) & wbMult(2486 downto 2484)) + (wbMult(2489) & wbMult(2489 downto 2487));
      v.Lvl1(1663 downto 1660) := (wbMult(2492) & wbMult(2492 downto 2490)) + (wbMult(2495) & wbMult(2495 downto 2493));
      v.Lvl1(1667 downto 1664) := (wbMult(2498) & wbMult(2498 downto 2496)) + (wbMult(2501) & wbMult(2501 downto 2499));
      v.Lvl1(1671 downto 1668) := (wbMult(2504) & wbMult(2504 downto 2502)) + (wbMult(2507) & wbMult(2507 downto 2505));
      v.Lvl1(1675 downto 1672) := (wbMult(2510) & wbMult(2510 downto 2508)) + (wbMult(2513) & wbMult(2513 downto 2511));
      v.Lvl1(1679 downto 1676) := (wbMult(2516) & wbMult(2516 downto 2514)) + (wbMult(2519) & wbMult(2519 downto 2517));
      v.Lvl1(1683 downto 1680) := (wbMult(2522) & wbMult(2522 downto 2520)) + (wbMult(2525) & wbMult(2525 downto 2523));
      v.Lvl1(1687 downto 1684) := (wbMult(2528) & wbMult(2528 downto 2526)) + (wbMult(2531) & wbMult(2531 downto 2529));
      v.Lvl1(1691 downto 1688) := (wbMult(2534) & wbMult(2534 downto 2532)) + (wbMult(2537) & wbMult(2537 downto 2535));
      v.Lvl1(1695 downto 1692) := (wbMult(2540) & wbMult(2540 downto 2538)) + (wbMult(2543) & wbMult(2543 downto 2541));
      v.Lvl1(1699 downto 1696) := (wbMult(2546) & wbMult(2546 downto 2544)) + (wbMult(2549) & wbMult(2549 downto 2547));
      v.Lvl1(1703 downto 1700) := (wbMult(2552) & wbMult(2552 downto 2550)) + (wbMult(2555) & wbMult(2555 downto 2553));
      v.Lvl1(1707 downto 1704) := (wbMult(2558) & wbMult(2558 downto 2556)) + (wbMult(2561) & wbMult(2561 downto 2559));
      v.Lvl1(1711 downto 1708) := (wbMult(2564) & wbMult(2564 downto 2562)) + (wbMult(2567) & wbMult(2567 downto 2565));
      v.Lvl1(1715 downto 1712) := (wbMult(2570) & wbMult(2570 downto 2568)) + (wbMult(2573) & wbMult(2573 downto 2571));
      v.Lvl1(1719 downto 1716) := (wbMult(2576) & wbMult(2576 downto 2574)) + (wbMult(2579) & wbMult(2579 downto 2577));
      v.Lvl1(1723 downto 1720) := (wbMult(2582) & wbMult(2582 downto 2580)) + (wbMult(2585) & wbMult(2585 downto 2583));
      v.Lvl1(1727 downto 1724) := (wbMult(2588) & wbMult(2588 downto 2586)) + (wbMult(2591) & wbMult(2591 downto 2589));
      v.Lvl1(1731 downto 1728) := (wbMult(2594) & wbMult(2594 downto 2592)) + (wbMult(2597) & wbMult(2597 downto 2595));
      v.Lvl1(1735 downto 1732) := (wbMult(2600) & wbMult(2600 downto 2598)) + (wbMult(2603) & wbMult(2603 downto 2601));
      v.Lvl1(1739 downto 1736) := (wbMult(2606) & wbMult(2606 downto 2604)) + (wbMult(2609) & wbMult(2609 downto 2607));
      v.Lvl1(1743 downto 1740) := (wbMult(2612) & wbMult(2612 downto 2610)) + (wbMult(2615) & wbMult(2615 downto 2613));
      v.Lvl1(1747 downto 1744) := (wbMult(2618) & wbMult(2618 downto 2616)) + (wbMult(2621) & wbMult(2621 downto 2619));
      v.Lvl1(1751 downto 1748) := (wbMult(2624) & wbMult(2624 downto 2622)) + (wbMult(2627) & wbMult(2627 downto 2625));
      v.Lvl1(1755 downto 1752) := (wbMult(2630) & wbMult(2630 downto 2628)) + (wbMult(2633) & wbMult(2633 downto 2631));
      v.Lvl1(1759 downto 1756) := (wbMult(2636) & wbMult(2636 downto 2634)) + (wbMult(2639) & wbMult(2639 downto 2637));
      v.Lvl1(1763 downto 1760) := (wbMult(2642) & wbMult(2642 downto 2640)) + (wbMult(2645) & wbMult(2645 downto 2643));
      v.Lvl1(1767 downto 1764) := (wbMult(2648) & wbMult(2648 downto 2646)) + (wbMult(2651) & wbMult(2651 downto 2649));
      v.Lvl1(1771 downto 1768) := (wbMult(2654) & wbMult(2654 downto 2652)) + (wbMult(2657) & wbMult(2657 downto 2655));
      v.Lvl1(1775 downto 1772) := (wbMult(2660) & wbMult(2660 downto 2658)) + (wbMult(2663) & wbMult(2663 downto 2661));
      v.Lvl1(1779 downto 1776) := (wbMult(2666) & wbMult(2666 downto 2664)) + (wbMult(2669) & wbMult(2669 downto 2667));
      v.Lvl1(1783 downto 1780) := (wbMult(2672) & wbMult(2672 downto 2670)) + (wbMult(2675) & wbMult(2675 downto 2673));
      v.Lvl1(1787 downto 1784) := (wbMult(2678) & wbMult(2678 downto 2676)) + (wbMult(2681) & wbMult(2681 downto 2679));
      v.Lvl1(1791 downto 1788) := (wbMult(2684) & wbMult(2684 downto 2682)) + (wbMult(2687) & wbMult(2687 downto 2685));
      v.Lvl1(1795 downto 1792) := (wbMult(2690) & wbMult(2690 downto 2688)) + (wbMult(2693) & wbMult(2693 downto 2691));
      v.Lvl1(1799 downto 1796) := (wbMult(2696) & wbMult(2696 downto 2694)) + (wbMult(2699) & wbMult(2699 downto 2697));
      v.Lvl1(1803 downto 1800) := (wbMult(2702) & wbMult(2702 downto 2700)) + (wbMult(2705) & wbMult(2705 downto 2703));
      v.Lvl1(1807 downto 1804) := (wbMult(2708) & wbMult(2708 downto 2706)) + (wbMult(2711) & wbMult(2711 downto 2709));
      v.Lvl1(1811 downto 1808) := (wbMult(2714) & wbMult(2714 downto 2712)) + (wbMult(2717) & wbMult(2717 downto 2715));
      v.Lvl1(1815 downto 1812) := (wbMult(2720) & wbMult(2720 downto 2718)) + (wbMult(2723) & wbMult(2723 downto 2721));
      v.Lvl1(1819 downto 1816) := (wbMult(2726) & wbMult(2726 downto 2724)) + (wbMult(2729) & wbMult(2729 downto 2727));
      v.Lvl1(1823 downto 1820) := (wbMult(2732) & wbMult(2732 downto 2730)) + (wbMult(2735) & wbMult(2735 downto 2733));
      v.Lvl1(1827 downto 1824) := (wbMult(2738) & wbMult(2738 downto 2736)) + (wbMult(2741) & wbMult(2741 downto 2739));
      v.Lvl1(1831 downto 1828) := (wbMult(2744) & wbMult(2744 downto 2742)) + (wbMult(2747) & wbMult(2747 downto 2745));
      v.Lvl1(1835 downto 1832) := (wbMult(2750) & wbMult(2750 downto 2748)) + (wbMult(2753) & wbMult(2753 downto 2751));
      v.Lvl1(1839 downto 1836) := (wbMult(2756) & wbMult(2756 downto 2754)) + (wbMult(2759) & wbMult(2759 downto 2757));
      v.Lvl1(1843 downto 1840) := (wbMult(2762) & wbMult(2762 downto 2760)) + (wbMult(2765) & wbMult(2765 downto 2763));
      v.Lvl1(1847 downto 1844) := (wbMult(2768) & wbMult(2768 downto 2766)) + (wbMult(2771) & wbMult(2771 downto 2769));
      v.Lvl1(1851 downto 1848) := (wbMult(2774) & wbMult(2774 downto 2772)) + (wbMult(2777) & wbMult(2777 downto 2775));
      v.Lvl1(1855 downto 1852) := (wbMult(2780) & wbMult(2780 downto 2778)) + (wbMult(2783) & wbMult(2783 downto 2781));
      v.Lvl1(1859 downto 1856) := (wbMult(2786) & wbMult(2786 downto 2784)) + (wbMult(2789) & wbMult(2789 downto 2787));
      v.Lvl1(1863 downto 1860) := (wbMult(2792) & wbMult(2792 downto 2790)) + (wbMult(2795) & wbMult(2795 downto 2793));
      v.Lvl1(1867 downto 1864) := (wbMult(2798) & wbMult(2798 downto 2796)) + (wbMult(2801) & wbMult(2801 downto 2799));
      v.Lvl1(1871 downto 1868) := (wbMult(2804) & wbMult(2804 downto 2802)) + (wbMult(2807) & wbMult(2807 downto 2805));
      v.Lvl1(1875 downto 1872) := (wbMult(2810) & wbMult(2810 downto 2808)) + (wbMult(2813) & wbMult(2813 downto 2811));
      v.Lvl1(1879 downto 1876) := (wbMult(2816) & wbMult(2816 downto 2814)) + (wbMult(2819) & wbMult(2819 downto 2817));
      v.Lvl1(1883 downto 1880) := (wbMult(2822) & wbMult(2822 downto 2820)) + (wbMult(2825) & wbMult(2825 downto 2823));
      v.Lvl1(1887 downto 1884) := (wbMult(2828) & wbMult(2828 downto 2826)) + (wbMult(2831) & wbMult(2831 downto 2829));
      v.Lvl1(1891 downto 1888) := (wbMult(2834) & wbMult(2834 downto 2832)) + (wbMult(2837) & wbMult(2837 downto 2835));
      v.Lvl1(1895 downto 1892) := (wbMult(2840) & wbMult(2840 downto 2838)) + (wbMult(2843) & wbMult(2843 downto 2841));
      v.Lvl1(1899 downto 1896) := (wbMult(2846) & wbMult(2846 downto 2844)) + (wbMult(2849) & wbMult(2849 downto 2847));
      v.Lvl1(1903 downto 1900) := (wbMult(2852) & wbMult(2852 downto 2850)) + (wbMult(2855) & wbMult(2855 downto 2853));
      v.Lvl1(1907 downto 1904) := (wbMult(2858) & wbMult(2858 downto 2856)) + (wbMult(2861) & wbMult(2861 downto 2859));
      v.Lvl1(1911 downto 1908) := (wbMult(2864) & wbMult(2864 downto 2862)) + (wbMult(2867) & wbMult(2867 downto 2865));
      v.Lvl1(1915 downto 1912) := (wbMult(2870) & wbMult(2870 downto 2868)) + (wbMult(2873) & wbMult(2873 downto 2871));
      v.Lvl1(1919 downto 1916) := (wbMult(2876) & wbMult(2876 downto 2874)) + (wbMult(2879) & wbMult(2879 downto 2877));
      v.Lvl1(1923 downto 1920) := (wbMult(2882) & wbMult(2882 downto 2880)) + (wbMult(2885) & wbMult(2885 downto 2883));
      v.Lvl1(1927 downto 1924) := (wbMult(2888) & wbMult(2888 downto 2886)) + (wbMult(2891) & wbMult(2891 downto 2889));
      v.Lvl1(1931 downto 1928) := (wbMult(2894) & wbMult(2894 downto 2892)) + (wbMult(2897) & wbMult(2897 downto 2895));
      v.Lvl1(1935 downto 1932) := (wbMult(2900) & wbMult(2900 downto 2898)) + (wbMult(2903) & wbMult(2903 downto 2901));
      v.Lvl1(1939 downto 1936) := (wbMult(2906) & wbMult(2906 downto 2904)) + (wbMult(2909) & wbMult(2909 downto 2907));
      v.Lvl1(1943 downto 1940) := (wbMult(2912) & wbMult(2912 downto 2910)) + (wbMult(2915) & wbMult(2915 downto 2913));
      v.Lvl1(1947 downto 1944) := (wbMult(2918) & wbMult(2918 downto 2916)) + (wbMult(2921) & wbMult(2921 downto 2919));
      v.Lvl1(1951 downto 1948) := (wbMult(2924) & wbMult(2924 downto 2922)) + (wbMult(2927) & wbMult(2927 downto 2925));
      v.Lvl1(1955 downto 1952) := (wbMult(2930) & wbMult(2930 downto 2928)) + (wbMult(2933) & wbMult(2933 downto 2931));
      v.Lvl1(1959 downto 1956) := (wbMult(2936) & wbMult(2936 downto 2934)) + (wbMult(2939) & wbMult(2939 downto 2937));
      v.Lvl1(1963 downto 1960) := (wbMult(2942) & wbMult(2942 downto 2940)) + (wbMult(2945) & wbMult(2945 downto 2943));
      v.Lvl1(1967 downto 1964) := (wbMult(2948) & wbMult(2948 downto 2946)) + (wbMult(2951) & wbMult(2951 downto 2949));
      v.Lvl1(1971 downto 1968) := (wbMult(2954) & wbMult(2954 downto 2952)) + (wbMult(2957) & wbMult(2957 downto 2955));
      v.Lvl1(1975 downto 1972) := (wbMult(2960) & wbMult(2960 downto 2958)) + (wbMult(2963) & wbMult(2963 downto 2961));
      v.Lvl1(1979 downto 1976) := (wbMult(2966) & wbMult(2966 downto 2964)) + (wbMult(2969) & wbMult(2969 downto 2967));
      v.Lvl1(1983 downto 1980) := (wbMult(2972) & wbMult(2972 downto 2970)) + (wbMult(2975) & wbMult(2975 downto 2973));
      v.Lvl1(1987 downto 1984) := (wbMult(2978) & wbMult(2978 downto 2976)) + (wbMult(2981) & wbMult(2981 downto 2979));
      v.Lvl1(1991 downto 1988) := (wbMult(2984) & wbMult(2984 downto 2982)) + (wbMult(2987) & wbMult(2987 downto 2985));
      v.Lvl1(1995 downto 1992) := (wbMult(2990) & wbMult(2990 downto 2988)) + (wbMult(2993) & wbMult(2993 downto 2991));
      v.Lvl1(1999 downto 1996) := (wbMult(2996) & wbMult(2996 downto 2994)) + (wbMult(2999) & wbMult(2999 downto 2997));
      v.Lvl1(2003 downto 2000) := (wbMult(3002) & wbMult(3002 downto 3000)) + (wbMult(3005) & wbMult(3005 downto 3003));
      v.Lvl1(2007 downto 2004) := (wbMult(3008) & wbMult(3008 downto 3006)) + (wbMult(3011) & wbMult(3011 downto 3009));
      v.Lvl1(2011 downto 2008) := (wbMult(3014) & wbMult(3014 downto 3012)) + (wbMult(3017) & wbMult(3017 downto 3015));
      v.Lvl1(2015 downto 2012) := (wbMult(3020) & wbMult(3020 downto 3018)) + (wbMult(3023) & wbMult(3023 downto 3021));
      v.Lvl1(2019 downto 2016) := (wbMult(3026) & wbMult(3026 downto 3024)) + (wbMult(3029) & wbMult(3029 downto 3027));
      v.Lvl1(2023 downto 2020) := (wbMult(3032) & wbMult(3032 downto 3030)) + (wbMult(3035) & wbMult(3035 downto 3033));
      v.Lvl1(2027 downto 2024) := (wbMult(3038) & wbMult(3038 downto 3036)) + (wbMult(3041) & wbMult(3041 downto 3039));
      v.Lvl1(2031 downto 2028) := (wbMult(3044) & wbMult(3044 downto 3042)) + (wbMult(3047) & wbMult(3047 downto 3045));
      v.Lvl1(2035 downto 2032) := (wbMult(3050) & wbMult(3050 downto 3048)) + (wbMult(3053) & wbMult(3053 downto 3051));
      v.Lvl1(2039 downto 2036) := (wbMult(3056) & wbMult(3056 downto 3054)) + (wbMult(3059) & wbMult(3059 downto 3057));
      v.Lvl1(2043 downto 2040) := (wbMult(3062) & wbMult(3062 downto 3060)) + (wbMult(3065) & wbMult(3065 downto 3063));
      v.Lvl1(2047 downto 2044) := (wbMult(3068) & wbMult(3068 downto 3066)) + (wbMult(3071) & wbMult(3071 downto 3069));
    --end if;

    if i_nrst = '0' then
      v.Lvl1 := (others => '0');
    end if;
    
    rin <= v;
  end process;
  

  o_lvl1 <= r.Lvl1;


  regs : process(i_clk)
  begin 
    if rising_edge(i_clk) then 
      r <= rin;
    end if;
  end process;

end; 

