//--------------------------------------------------------------------------
//! @author     Sergey Khabarov
//! @brief      Virtual simple output buffer.
//--------------------------------------------------------------------------

module obuf_tech (
    output logic o,
    input i
); 
 
    assign o = i;

endmodule
