//--------------------------------------------------------------------------
//! @author     Sergey Khabarov
//! @brief      Virtual simple input buffer.
//----------------------------------------------------------------------------

module ibuf_tech(
    output logic o,
    input i
);

   assign o = i;
   
endmodule
