//--------------------------------------------------------------------------
//! @author     Sergey Khabarov
//! @brief      Virtual clock buffered output.
//----------------------------------------------------------------------------

module ibufg_tech (
    output logic o,
    input i
);

    assign o = i;

endmodule
