module Htif(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_csr,
    output io_cpu_0_reset,
    output io_cpu_0_id,
    input  io_cpu_0_csr_req_ready,
    output io_cpu_0_csr_req_valid,
    output io_cpu_0_csr_req_bits_rw,
    output[11:0] io_cpu_0_csr_req_bits_addr,
    output[63:0] io_cpu_0_csr_req_bits_data,
    output io_cpu_0_csr_resp_ready,
    input  io_cpu_0_csr_resp_valid,
    input [63:0] io_cpu_0_csr_resp_bits,
    output io_cpu_0_ipi_req_ready,
    input  io_cpu_0_ipi_req_valid,
    input  io_cpu_0_ipi_req_bits,
    input  io_cpu_0_ipi_rep_ready,
    output io_cpu_0_ipi_rep_valid,
    //output io_cpu_0_ipi_rep_bits
    input  io_cpu_0_debug_stats_csr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[1:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_scr_req_ready,
    output io_scr_req_valid,
    output io_scr_req_bits_rw,
    output[5:0] io_scr_req_bits_addr,
    output[63:0] io_scr_req_bits_data,
    output io_scr_resp_ready,
    input  io_scr_resp_valid,
    input [63:0] io_scr_resp_bits
);

  wire[63:0] csr_wdata;
  reg [63:0] packet_ram [7:0];
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire T3;
  reg [2:0] state;
  wire[2:0] T215;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire T18;
  wire T19;
  wire[3:0] rx_cmd;
  reg [3:0] cmd;
  wire[3:0] T20;
  wire T21;
  wire T22;
  reg [14:0] rx_count;
  wire[14:0] T216;
  wire[14:0] T23;
  wire[14:0] T24;
  wire[14:0] T25;
  wire T26;
  wire T27;
  wire[12:0] T217;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T28;
  wire[11:0] T29;
  wire[63:0] rx_shifter_in;
  wire[47:0] T30;
  reg [63:0] rx_shifter;
  wire[63:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire nack;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire bad_mem_packet;
  wire T44;
  wire[2:0] T45;
  reg [39:0] addr;
  wire[39:0] T46;
  wire[39:0] T47;
  wire[39:0] T48;
  wire[39:0] T49;
  wire[39:0] T50;
  wire[39:0] T51;
  wire T52;
  wire[2:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire[12:0] tx_word_count;
  reg [14:0] tx_count;
  wire[14:0] T218;
  wire[14:0] T57;
  wire[14:0] T58;
  wire[14:0] T59;
  wire T60;
  wire T61;
  wire[3:0] next_cmd;
  wire T62;
  wire[12:0] rx_word_count;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire rx_done;
  wire T67;
  wire T68;
  wire T69;
  wire[2:0] T70;
  wire T71;
  wire[12:0] T219;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire rx_word_done;
  wire T76;
  wire[1:0] T77;
  wire T78;
  wire T79;
  wire cnt_done;
  wire T80;
  reg [1:0] cnt;
  wire[1:0] T220;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  reg [8:0] pos;
  wire[8:0] T94;
  wire[8:0] T95;
  wire[8:0] T96;
  wire[8:0] T97;
  wire[8:0] T98;
  wire[8:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[2:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[2:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire tx_done;
  wire T114;
  wire T115;
  wire T116;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T117;
  wire T118;
  wire T119;
  wire[12:0] T221;
  wire T120;
  wire T121;
  wire[1:0] tx_subword_count;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire[11:0] csr_addr;
  wire T126;
  wire T127;
  wire[1:0] csr_coreid;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[63:0] T135;
  wire[63:0] T136;
  wire T137;
  wire T138;
  wire[2:0] T139;
  wire[63:0] T140;
  wire T141;
  wire[2:0] T142;
  wire[2:0] T143;
  wire[5:0] T144;
  wire[5:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[127:0] T150;
  wire[127:0] T151;
  wire[127:0] T152;
  wire[127:0] mem_req_data;
  wire[63:0] T153;
  wire[2:0] T154;
  wire[63:0] T155;
  wire[2:0] T156;
  wire T157;
  wire[16:0] T158;
  wire[16:0] T159;
  wire[16:0] T160;
  wire[16:0] T161;
  wire[15:0] T162;
  wire[2:0] T163;
  wire[2:0] T164;
  wire[2:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[1:0] T171;
  wire[1:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire[25:0] T175;
  wire[25:0] T176;
  wire[25:0] T222;
  wire[36:0] init_addr;
  wire[39:0] T177;
  wire[25:0] T178;
  wire[25:0] T223;
  wire T179;
  wire T180;
  wire T181;
  reg  R182;
  wire T224;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  R192;
  wire T225;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[15:0] T226;
  wire[63:0] T197;
  wire[5:0] T198;
  wire[1:0] T199;
  wire[63:0] tx_data;
  wire[63:0] T200;
  wire[63:0] T201;
  reg [63:0] csrReadData;
  wire[63:0] T202;
  wire[63:0] T203;
  wire[63:0] T204;
  wire[63:0] T227;
  wire T205;
  wire T206;
  wire T207;
  wire[63:0] tx_header;
  wire[15:0] T208;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T209;
  reg [7:0] seqno;
  wire[7:0] T210;
  wire[7:0] T211;
  wire T212;
  wire T213;
  wire T214;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    state = {1{$random}};
    cmd = {1{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    rx_shifter = {2{$random}};
    addr = {2{$random}};
    tx_count = {1{$random}};
    cnt = {1{$random}};
    pos = {1{$random}};
    R182 = {1{$random}};
    R192 = {1{$random}};
    csrReadData = {2{$random}};
    seqno = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_cpu_0_ipi_rep_bits = {1{$random}};
  assign io_cpu_0_id = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_scr_resp_ready = 1'h1;
  assign io_scr_req_bits_data = csr_wdata;
  assign csr_wdata = packet_ram[3'h0];
  assign T1 = io_mem_grant_bits_data[7'h7f:7'h40];
  assign T2 = T3 & io_mem_grant_valid;
  assign T3 = state == 3'h5;
  assign T215 = reset ? 3'h0 : T4;
  assign T4 = T132 ? 3'h7 : T5;
  assign T5 = T131 ? 3'h2 : T6;
  assign T6 = T129 ? 3'h7 : T7;
  assign T7 = T124 ? 3'h7 : T8;
  assign T8 = T123 ? 3'h2 : T9;
  assign T9 = T113 ? T109 : T10;
  assign T10 = T107 ? T103 : T11;
  assign T11 = T101 ? T91 : T12;
  assign T12 = T89 ? 3'h5 : T13;
  assign T13 = T79 ? 3'h6 : T14;
  assign T14 = T66 ? T15 : state;
  assign T15 = T65 ? 3'h3 : T16;
  assign T16 = T64 ? 3'h4 : T17;
  assign T17 = T18 ? 3'h1 : 3'h7;
  assign T18 = T63 | T19;
  assign T19 = rx_cmd == 4'h3;
  assign rx_cmd = T62 ? next_cmd : cmd;
  assign T20 = T21 ? next_cmd : cmd;
  assign T21 = T61 & T22;
  assign T22 = rx_count == 15'h3;
  assign T216 = reset ? 15'h0 : T23;
  assign T23 = T26 ? 15'h0 : T24;
  assign T24 = T61 ? T25 : rx_count;
  assign T25 = rx_count + 15'h1;
  assign T26 = T113 & T27;
  assign T27 = tx_word_count == T217;
  assign T217 = {1'h0, tx_size};
  assign tx_size = T32 ? size : 12'h0;
  assign T28 = T21 ? T29 : size;
  assign T29 = rx_shifter_in[4'hf:3'h4];
  assign rx_shifter_in = {io_host_in_bits, T30};
  assign T30 = rx_shifter[6'h3f:5'h10];
  assign T31 = T61 ? rx_shifter_in : rx_shifter;
  assign T32 = T38 & T33;
  assign T33 = T35 | T34;
  assign T34 = cmd == 4'h3;
  assign T35 = T37 | T36;
  assign T36 = cmd == 4'h2;
  assign T37 = cmd == 4'h0;
  assign T38 = nack ^ 1'h1;
  assign nack = T54 ? bad_mem_packet : T39;
  assign T39 = T41 ? T40 : 1'h1;
  assign T40 = size != 12'h1;
  assign T41 = T43 | T42;
  assign T42 = cmd == 4'h3;
  assign T43 = cmd == 4'h2;
  assign bad_mem_packet = T52 | T44;
  assign T44 = T45 != 3'h0;
  assign T45 = addr[2'h2:1'h0];
  assign T46 = T107 ? T51 : T47;
  assign T47 = T101 ? T50 : T48;
  assign T48 = T21 ? T49 : addr;
  assign T49 = rx_shifter_in[6'h3f:5'h18];
  assign T50 = addr + 40'h8;
  assign T51 = addr + 40'h8;
  assign T52 = T53 != 3'h0;
  assign T53 = size[2'h2:1'h0];
  assign T54 = T56 | T55;
  assign T55 = cmd == 4'h1;
  assign T56 = cmd == 4'h0;
  assign tx_word_count = tx_count[4'he:2'h2];
  assign T218 = reset ? 15'h0 : T57;
  assign T57 = T26 ? 15'h0 : T58;
  assign T58 = T60 ? T59 : tx_count;
  assign T59 = tx_count + 15'h1;
  assign T60 = io_host_out_valid & io_host_out_ready;
  assign T61 = io_host_in_valid & io_host_in_ready;
  assign next_cmd = rx_shifter_in[2'h3:1'h0];
  assign T62 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T63 = rx_cmd == 4'h2;
  assign T64 = rx_cmd == 4'h1;
  assign T65 = rx_cmd == 4'h0;
  assign T66 = T78 & rx_done;
  assign rx_done = rx_word_done & T67;
  assign T67 = T75 ? T72 : T68;
  assign T68 = T71 | T69;
  assign T69 = T70 == 3'h0;
  assign T70 = rx_word_count[2'h2:1'h0];
  assign T71 = rx_word_count == T219;
  assign T219 = {1'h0, size};
  assign T72 = T74 & T73;
  assign T73 = next_cmd != 4'h3;
  assign T74 = next_cmd != 4'h1;
  assign T75 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T76;
  assign T76 = T77 == 2'h3;
  assign T77 = rx_count[1'h1:1'h0];
  assign T78 = state == 3'h0;
  assign T79 = T88 & cnt_done;
  assign cnt_done = T83 & T80;
  assign T80 = cnt == 2'h3;
  assign T220 = reset ? 2'h0 : T81;
  assign T81 = T83 ? T82 : cnt;
  assign T82 = cnt + 2'h1;
  assign T83 = T86 | T84;
  assign T84 = T85 & io_mem_grant_valid;
  assign T85 = state == 3'h5;
  assign T86 = T87 & io_mem_acquire_ready;
  assign T87 = state == 3'h4;
  assign T88 = state == 3'h4;
  assign T89 = T90 & io_mem_acquire_ready;
  assign T90 = state == 3'h3;
  assign T91 = T92 ? 3'h7 : 3'h0;
  assign T92 = T100 | T93;
  assign T93 = pos == 9'h1;
  assign T94 = T107 ? T99 : T95;
  assign T95 = T101 ? T98 : T96;
  assign T96 = T21 ? T97 : pos;
  assign T97 = rx_shifter_in[4'hf:3'h7];
  assign T98 = pos - 9'h1;
  assign T99 = pos - 9'h1;
  assign T100 = cmd == 4'h0;
  assign T101 = T102 & io_mem_grant_valid;
  assign T102 = state == 3'h6;
  assign T103 = T104 ? 3'h7 : 3'h0;
  assign T104 = T106 | T105;
  assign T105 = pos == 9'h1;
  assign T106 = cmd == 4'h0;
  assign T107 = T108 & cnt_done;
  assign T108 = state == 3'h5;
  assign T109 = T110 ? 3'h3 : 3'h0;
  assign T110 = T112 & T111;
  assign T111 = pos != 9'h0;
  assign T112 = cmd == 4'h0;
  assign T113 = T122 & tx_done;
  assign tx_done = T120 & T114;
  assign T114 = T119 | T115;
  assign T115 = T118 & T116;
  assign T116 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T117 - 3'h1;
  assign T117 = tx_word_count[2'h2:1'h0];
  assign T118 = 13'h0 < tx_word_count;
  assign T119 = tx_word_count == T221;
  assign T221 = {1'h0, tx_size};
  assign T120 = io_host_out_ready & T121;
  assign T121 = tx_subword_count == 2'h3;
  assign tx_subword_count = tx_count[1'h1:1'h0];
  assign T122 = state == 3'h7;
  assign T123 = io_cpu_0_csr_req_ready & io_cpu_0_csr_req_valid;
  assign T124 = T126 & T125;
  assign T125 = csr_addr == 12'h782;
  assign csr_addr = addr[4'hb:1'h0];
  assign T126 = T128 & T127;
  assign T127 = csr_coreid == 2'h0;
  assign csr_coreid = addr[5'h15:5'h14];
  assign T128 = state == 3'h1;
  assign T129 = T130 & io_cpu_0_csr_resp_valid;
  assign T130 = state == 3'h2;
  assign T131 = io_scr_req_ready & io_scr_req_valid;
  assign T132 = T133 & io_scr_resp_valid;
  assign T133 = state == 3'h2;
  assign T134 = {io_mem_grant_bits_addr_beat, 1'h1};
  assign T136 = io_mem_grant_bits_data[6'h3f:1'h0];
  assign T137 = T138 & io_mem_grant_valid;
  assign T138 = state == 3'h5;
  assign T139 = {io_mem_grant_bits_addr_beat, 1'h0};
  assign T141 = rx_word_done & io_host_in_ready;
  assign T142 = T143 - 3'h1;
  assign T143 = rx_word_count[2'h2:1'h0];
  assign io_scr_req_bits_addr = T144;
  assign T144 = T145;
  assign T145 = addr[3'h5:1'h0];
  assign io_scr_req_bits_rw = T146;
  assign T146 = cmd == 4'h3;
  assign io_scr_req_valid = T147;
  assign T147 = T149 & T148;
  assign T148 = csr_coreid == 2'h3;
  assign T149 = state == 3'h1;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_data = T150;
  assign T150 = T157 ? T152 : T151;
  assign T151 = 128'h0;
  assign T152 = mem_req_data;
  assign mem_req_data = {T155, T153};
  assign T153 = packet_ram[T154];
  assign T154 = {cnt, 1'h0};
  assign T155 = packet_ram[T156];
  assign T156 = {cnt, 1'h1};
  assign T157 = cmd == 4'h1;
  assign io_mem_acquire_bits_union = T158;
  assign T158 = T157 ? T160 : T159;
  assign T159 = 17'h1c1;
  assign T160 = T161;
  assign T161 = {T162, 1'h1};
  assign T162 = 16'hffff;
  assign io_mem_acquire_bits_a_type = T163;
  assign T163 = T157 ? T165 : T164;
  assign T164 = 3'h1;
  assign T165 = 3'h3;
  assign io_mem_acquire_bits_is_builtin_type = T166;
  assign T166 = T157 ? T168 : T167;
  assign T167 = 1'h1;
  assign T168 = 1'h1;
  assign io_mem_acquire_bits_addr_beat = T169;
  assign T169 = T157 ? T171 : T170;
  assign T170 = 2'h0;
  assign T171 = cnt;
  assign io_mem_acquire_bits_client_xact_id = T172;
  assign T172 = T157 ? T174 : T173;
  assign T173 = 2'h0;
  assign T174 = 2'h0;
  assign io_mem_acquire_bits_addr_block = T175;
  assign T175 = T157 ? T178 : T176;
  assign T176 = T222;
  assign T222 = init_addr[5'h19:1'h0];
  assign init_addr = T177 >> 2'h3;
  assign T177 = addr;
  assign T178 = T223;
  assign T223 = init_addr[5'h19:1'h0];
  assign io_mem_acquire_valid = T179;
  assign T179 = T181 | T180;
  assign T180 = state == 3'h4;
  assign T181 = state == 3'h3;
  assign io_cpu_0_ipi_rep_valid = R182;
  assign T224 = reset ? 1'h0 : T183;
  assign T183 = T185 ? 1'h1 : T184;
  assign T184 = io_cpu_0_ipi_rep_ready ? 1'h0 : R182;
  assign T185 = io_cpu_0_ipi_req_valid & T186;
  assign T186 = io_cpu_0_ipi_req_bits == 1'h0;
  assign io_cpu_0_ipi_req_ready = 1'h1;
  assign io_cpu_0_csr_resp_ready = 1'h1;
  assign io_cpu_0_csr_req_bits_data = csr_wdata;
  assign io_cpu_0_csr_req_bits_addr = csr_addr;
  assign io_cpu_0_csr_req_bits_rw = T187;
  assign T187 = cmd == 4'h3;
  assign io_cpu_0_csr_req_valid = T188;
  assign T188 = T190 & T189;
  assign T189 = csr_addr != 12'h782;
  assign T190 = T191 & T127;
  assign T191 = state == 3'h1;
  assign io_cpu_0_reset = R192;
  assign T225 = reset ? 1'h1 : T193;
  assign T193 = T195 ? T194 : R192;
  assign T194 = csr_wdata[1'h0:1'h0];
  assign T195 = T124 & T196;
  assign T196 = cmd == 4'h3;
  assign io_host_debug_stats_csr = io_cpu_0_debug_stats_csr;
  assign io_host_out_bits = T226;
  assign T226 = T197[4'hf:1'h0];
  assign T197 = tx_data >> T198;
  assign T198 = {T199, 4'h0};
  assign T199 = tx_count[1'h1:1'h0];
  assign tx_data = T212 ? tx_header : T200;
  assign T200 = T205 ? csrReadData : T201;
  assign T201 = packet_ram[packet_ram_raddr];
  assign T202 = T132 ? io_scr_resp_bits : T203;
  assign T203 = T129 ? io_cpu_0_csr_resp_bits : T204;
  assign T204 = T124 ? T227 : csrReadData;
  assign T227 = {63'h0, R192};
  assign T205 = T207 | T206;
  assign T206 = cmd == 4'h3;
  assign T207 = cmd == 4'h2;
  assign tx_header = {T209, T208};
  assign T208 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T209 = {addr, seqno};
  assign T210 = T21 ? T211 : seqno;
  assign T211 = rx_shifter_in[5'h17:5'h10];
  assign T212 = tx_word_count == 13'h0;
  assign io_host_out_valid = T213;
  assign T213 = state == 3'h7;
  assign io_host_in_ready = T214;
  assign T214 = state == 3'h0;

  always @(posedge clk) begin
    if (T2)
      packet_ram[T134] <= T1;
    if(reset) begin
      state <= 3'h0;
    end else if(T132) begin
      state <= 3'h7;
    end else if(T131) begin
      state <= 3'h2;
    end else if(T129) begin
      state <= 3'h7;
    end else if(T124) begin
      state <= 3'h7;
    end else if(T123) begin
      state <= 3'h2;
    end else if(T113) begin
      state <= T109;
    end else if(T107) begin
      state <= T103;
    end else if(T101) begin
      state <= T91;
    end else if(T89) begin
      state <= 3'h5;
    end else if(T79) begin
      state <= 3'h6;
    end else if(T66) begin
      state <= T15;
    end
    if(T21) begin
      cmd <= next_cmd;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T26) begin
      rx_count <= 15'h0;
    end else if(T61) begin
      rx_count <= T25;
    end
    if(T21) begin
      size <= T29;
    end
    if(T61) begin
      rx_shifter <= rx_shifter_in;
    end
    if(T107) begin
      addr <= T51;
    end else if(T101) begin
      addr <= T50;
    end else if(T21) begin
      addr <= T49;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T26) begin
      tx_count <= 15'h0;
    end else if(T60) begin
      tx_count <= T59;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T83) begin
      cnt <= T82;
    end
    if(T107) begin
      pos <= T99;
    end else if(T101) begin
      pos <= T98;
    end else if(T21) begin
      pos <= T97;
    end
    if (T137)
      packet_ram[T139] <= T136;
    if (T141)
      packet_ram[T142] <= rx_shifter_in;
    if(reset) begin
      R182 <= 1'h0;
    end else if(T185) begin
      R182 <= 1'h1;
    end else if(io_cpu_0_ipi_rep_ready) begin
      R182 <= 1'h0;
    end
    if(reset) begin
      R192 <= 1'h1;
    end else if(T195) begin
      R192 <= T194;
    end
    if(T132) begin
      csrReadData <= io_scr_resp_bits;
    end else if(T129) begin
      csrReadData <= io_cpu_0_csr_resp_bits;
    end else if(T124) begin
      csrReadData <= T227;
    end
    if(T21) begin
      seqno <= T211;
    end
  end
endmodule

module ClientTileLinkIOWrapper_0(
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [1:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[1:0] io_in_grant_bits_client_xact_id,
    output[3:0] io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[1:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [1:0] io_out_grant_bits_client_xact_id,
    input [3:0] io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [25:0] io_out_probe_bits_addr_block,
    input [1:0] io_out_probe_bits_p_type,
    input  io_out_release_ready,
    output io_out_release_valid
    //output[1:0] io_out_release_bits_addr_beat
    //output[25:0] io_out_release_bits_addr_block
    //output[1:0] io_out_release_bits_client_xact_id
    //output[2:0] io_out_release_bits_r_type
    //output io_out_release_bits_voluntary
    //output[127:0] io_out_release_bits_data
);



`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_out_release_bits_data = {4{$random}};
//  assign io_out_release_bits_voluntary = {1{$random}};
//  assign io_out_release_bits_r_type = {1{$random}};
//  assign io_out_release_bits_client_xact_id = {1{$random}};
//  assign io_out_release_bits_addr_block = {1{$random}};
//  assign io_out_release_bits_addr_beat = {1{$random}};
// synthesis translate_on
`endif
  assign io_out_release_valid = 1'h0;
  assign io_out_probe_ready = 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_in_grant_bits_data = io_out_grant_bits_data;
  assign io_in_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = io_out_acquire_ready;
endmodule

module FinishQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [3:0] io_enq_bits_fin_manager_xact_id,
    input [1:0] io_enq_bits_dst,
    input  io_deq_ready,
    output io_deq_valid,
    output[3:0] io_deq_bits_fin_manager_xact_id,
    output[1:0] io_deq_bits_dst,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T19;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T20;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T21;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[5:0] T11;
  reg [5:0] ram [1:0];
  wire[5:0] T12;
  wire[5:0] T13;
  wire[5:0] T14;
  wire[3:0] T15;
  wire T16;
  wire empty;
  wire T17;
  wire T18;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T19 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T20 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T21 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_dst = T10;
  assign T10 = T11[1'h1:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_fin_manager_xact_id, io_enq_bits_dst};
  assign io_deq_bits_fin_manager_xact_id = T15;
  assign T15 = T11[3'h5:2'h2];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module FinishUnit_0(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [1:0] io_grant_bits_header_src,
    input [1:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [1:0] io_grant_bits_payload_client_xact_id,
    input [3:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input [127:0] io_grant_bits_payload_data,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[1:0] io_refill_bits_client_xact_id,
    output[3:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    output[127:0] io_refill_bits_data,
    input  io_finish_ready,
    output io_finish_valid,
    output[1:0] io_finish_bits_header_src,
    output[1:0] io_finish_bits_header_dst,
    output[3:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[3:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T33;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[3:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[1:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T33 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 2'h0;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = io_grant_valid;
  assign io_grant_ready = T27;
  assign T27 = T28 & io_refill_ready;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_0(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [1:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[1:0] io_client_grant_bits_client_xact_id,
    output[3:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    output[127:0] io_client_grant_bits_data,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_addr_beat,
    input [25:0] io_client_release_bits_addr_block,
    input [1:0] io_client_release_bits_client_xact_id,
    input [2:0] io_client_release_bits_r_type,
    input  io_client_release_bits_voluntary,
    input [127:0] io_client_release_bits_data,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[1:0] io_network_acquire_bits_header_src,
    output[1:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[1:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [1:0] io_network_grant_bits_header_src,
    input [1:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [1:0] io_network_grant_bits_payload_client_xact_id,
    input [3:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[1:0] io_network_finish_bits_header_src,
    output[1:0] io_network_finish_bits_header_dst,
    output[3:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [1:0] io_network_probe_bits_header_src,
    input [1:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[1:0] io_network_release_bits_header_src,
    output[1:0] io_network_release_bits_header_dst,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[1:0] io_network_release_bits_payload_client_xact_id,
    output[2:0] io_network_release_bits_payload_r_type,
    output io_network_release_bits_payload_voluntary,
    output[127:0] io_network_release_bits_payload_data
);

  wire[127:0] rel_with_header_bits_payload_data;
  wire rel_with_header_bits_payload_voluntary;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire[1:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[1:0] rel_with_header_bits_header_dst;
  wire[1:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[1:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[1:0] acq_with_header_bits_header_dst;
  wire[1:0] acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[1:0] finisher_io_refill_bits_client_xact_id;
  wire[3:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_finish_valid;
  wire[1:0] finisher_io_finish_bits_header_src;
  wire[1:0] finisher_io_finish_bits_header_dst;
  wire[3:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 2'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 2'h0;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 2'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 2'h0;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_0 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [1:0] io_enq_bits_payload_addr_beat,
    input  io_enq_bits_payload_is_builtin_type,
    input [2:0] io_enq_bits_payload_a_type,
    input [16:0] io_enq_bits_payload_union,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[1:0] io_deq_bits_payload_addr_beat,
    output io_deq_bits_payload_is_builtin_type,
    output[2:0] io_deq_bits_payload_a_type,
    output[16:0] io_deq_bits_payload_union,
    output[127:0] io_deq_bits_payload_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T33;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T34;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T35;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[182:0] T11;
  reg [182:0] ram [1:0];
  wire[182:0] T12;
  wire[182:0] T13;
  wire[182:0] T14;
  wire[150:0] T15;
  wire[147:0] T16;
  wire[144:0] T17;
  wire[2:0] T18;
  wire[31:0] T19;
  wire[27:0] T20;
  wire[3:0] T21;
  wire[16:0] T22;
  wire[2:0] T23;
  wire T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[25:0] T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire T30;
  wire empty;
  wire T31;
  wire T32;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T33 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T34 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T35 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T19, T15};
  assign T15 = {T18, T16};
  assign T16 = {io_enq_bits_payload_a_type, T17};
  assign T17 = {io_enq_bits_payload_union, io_enq_bits_payload_data};
  assign T18 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_is_builtin_type};
  assign T19 = {T21, T20};
  assign T20 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_client_xact_id};
  assign T21 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_union = T22;
  assign T22 = T11[8'h90:8'h80];
  assign io_deq_bits_payload_a_type = T23;
  assign T23 = T11[8'h93:8'h91];
  assign io_deq_bits_payload_is_builtin_type = T24;
  assign T24 = T11[8'h94:8'h94];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'h96:8'h95];
  assign io_deq_bits_payload_client_xact_id = T26;
  assign T26 = T11[8'h98:8'h97];
  assign io_deq_bits_payload_addr_block = T27;
  assign T27 = T11[8'hb2:8'h99];
  assign io_deq_bits_header_dst = T28;
  assign T28 = T11[8'hb4:8'hb3];
  assign io_deq_bits_header_src = T29;
  assign T29 = T11[8'hb6:8'hb5];
  assign io_deq_valid = T30;
  assign T30 = empty ^ 1'h1;
  assign empty = ptr_match & T31;
  assign T31 = maybe_full ^ 1'h1;
  assign io_enq_ready = T32;
  assign T32 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_p_type,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T23;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T24;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T25;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[31:0] T11;
  reg [31:0] ram [1:0];
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[27:0] T15;
  wire[3:0] T16;
  wire[25:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire empty;
  wire T21;
  wire T22;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T23 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T24 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T25 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_p_type = T10;
  assign T10 = T11[1'h1:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T16, T15};
  assign T15 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_p_type};
  assign T16 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_addr_block = T17;
  assign T17 = T11[5'h1b:2'h2];
  assign io_deq_bits_header_dst = T18;
  assign T18 = T11[5'h1d:5'h1c];
  assign io_deq_bits_header_src = T19;
  assign T19 = T11[5'h1f:5'h1e];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_enq_bits_payload_voluntary,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_r_type,
    output io_deq_bits_payload_voluntary,
    output[127:0] io_deq_bits_payload_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T31;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T32;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[165:0] T11;
  reg [165:0] ram [1:0];
  wire[165:0] T12;
  wire[165:0] T13;
  wire[165:0] T14;
  wire[133:0] T15;
  wire[128:0] T16;
  wire[4:0] T17;
  wire[31:0] T18;
  wire[27:0] T19;
  wire[3:0] T20;
  wire T21;
  wire[2:0] T22;
  wire[1:0] T23;
  wire[25:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_voluntary, io_enq_bits_payload_data};
  assign T17 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_r_type};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_addr_block};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_voluntary = T21;
  assign T21 = T11[8'h80:8'h80];
  assign io_deq_bits_payload_r_type = T22;
  assign T22 = T11[8'h83:8'h81];
  assign io_deq_bits_payload_client_xact_id = T23;
  assign T23 = T11[8'h85:8'h84];
  assign io_deq_bits_payload_addr_block = T24;
  assign T24 = T11[8'h9f:8'h86];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'ha1:8'ha0];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[8'ha3:8'ha2];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[8'ha5:8'ha4];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [3:0] io_enq_bits_payload_manager_xact_id,
    input  io_enq_bits_payload_is_builtin_type,
    input [3:0] io_enq_bits_payload_g_type,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[3:0] io_deq_bits_payload_manager_xact_id,
    output io_deq_bits_payload_is_builtin_type,
    output[3:0] io_deq_bits_payload_g_type,
    output[127:0] io_deq_bits_payload_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T31;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T32;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[144:0] T11;
  reg [144:0] ram [1:0];
  wire[144:0] T12;
  wire[144:0] T13;
  wire[144:0] T14;
  wire[136:0] T15;
  wire[131:0] T16;
  wire[4:0] T17;
  wire[7:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire T22;
  wire[3:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_g_type, io_enq_bits_payload_data};
  assign T17 = {io_enq_bits_payload_manager_xact_id, io_enq_bits_payload_is_builtin_type};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_client_xact_id};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_g_type = T21;
  assign T21 = T11[8'h83:8'h80];
  assign io_deq_bits_payload_is_builtin_type = T22;
  assign T22 = T11[8'h84:8'h84];
  assign io_deq_bits_payload_manager_xact_id = T23;
  assign T23 = T11[8'h88:8'h85];
  assign io_deq_bits_payload_client_xact_id = T24;
  assign T24 = T11[8'h8a:8'h89];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'h8c:8'h8b];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[8'h8e:8'h8d];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[8'h90:8'h8f];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [3:0] io_enq_bits_payload_manager_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[3:0] io_deq_bits_payload_manager_xact_id,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[3:0] T10;
  wire[7:0] T11;
  reg [7:0] ram [1:0];
  wire[7:0] T12;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[5:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_manager_xact_id = T10;
  assign T10 = T11[2'h3:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_header_src, T15};
  assign T15 = {io_enq_bits_header_dst, io_enq_bits_payload_manager_xact_id};
  assign io_deq_bits_header_dst = T16;
  assign T16 = T11[3'h5:3'h4];
  assign io_deq_bits_header_src = T17;
  assign T17 = T11[3'h7:3'h6];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module TileLinkEnqueuer_0(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [1:0] io_client_acquire_bits_header_src,
    input [1:0] io_client_acquire_bits_header_dst,
    input [25:0] io_client_acquire_bits_payload_addr_block,
    input [1:0] io_client_acquire_bits_payload_client_xact_id,
    input [1:0] io_client_acquire_bits_payload_addr_beat,
    input  io_client_acquire_bits_payload_is_builtin_type,
    input [2:0] io_client_acquire_bits_payload_a_type,
    input [16:0] io_client_acquire_bits_payload_union,
    input [127:0] io_client_acquire_bits_payload_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_header_src,
    output[1:0] io_client_grant_bits_header_dst,
    output[1:0] io_client_grant_bits_payload_addr_beat,
    output[1:0] io_client_grant_bits_payload_client_xact_id,
    output[3:0] io_client_grant_bits_payload_manager_xact_id,
    output io_client_grant_bits_payload_is_builtin_type,
    output[3:0] io_client_grant_bits_payload_g_type,
    output[127:0] io_client_grant_bits_payload_data,
    output io_client_finish_ready,
    input  io_client_finish_valid,
    input [1:0] io_client_finish_bits_header_src,
    input [1:0] io_client_finish_bits_header_dst,
    input [3:0] io_client_finish_bits_payload_manager_xact_id,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[1:0] io_client_probe_bits_header_src,
    output[1:0] io_client_probe_bits_header_dst,
    output[25:0] io_client_probe_bits_payload_addr_block,
    output[1:0] io_client_probe_bits_payload_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_header_src,
    input [1:0] io_client_release_bits_header_dst,
    input [1:0] io_client_release_bits_payload_addr_beat,
    input [25:0] io_client_release_bits_payload_addr_block,
    input [1:0] io_client_release_bits_payload_client_xact_id,
    input [2:0] io_client_release_bits_payload_r_type,
    input  io_client_release_bits_payload_voluntary,
    input [127:0] io_client_release_bits_payload_data,
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[1:0] io_manager_acquire_bits_header_src,
    output[1:0] io_manager_acquire_bits_header_dst,
    output[25:0] io_manager_acquire_bits_payload_addr_block,
    output[1:0] io_manager_acquire_bits_payload_client_xact_id,
    output[1:0] io_manager_acquire_bits_payload_addr_beat,
    output io_manager_acquire_bits_payload_is_builtin_type,
    output[2:0] io_manager_acquire_bits_payload_a_type,
    output[16:0] io_manager_acquire_bits_payload_union,
    output[127:0] io_manager_acquire_bits_payload_data,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_header_src,
    input [1:0] io_manager_grant_bits_header_dst,
    input [1:0] io_manager_grant_bits_payload_addr_beat,
    input [1:0] io_manager_grant_bits_payload_client_xact_id,
    input [3:0] io_manager_grant_bits_payload_manager_xact_id,
    input  io_manager_grant_bits_payload_is_builtin_type,
    input [3:0] io_manager_grant_bits_payload_g_type,
    input [127:0] io_manager_grant_bits_payload_data,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[1:0] io_manager_finish_bits_header_src,
    output[1:0] io_manager_finish_bits_header_dst,
    output[3:0] io_manager_finish_bits_payload_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [1:0] io_manager_probe_bits_header_src,
    input [1:0] io_manager_probe_bits_header_dst,
    input [25:0] io_manager_probe_bits_payload_addr_block,
    input [1:0] io_manager_probe_bits_payload_p_type,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_header_src,
    output[1:0] io_manager_release_bits_header_dst,
    output[1:0] io_manager_release_bits_payload_addr_beat,
    output[25:0] io_manager_release_bits_payload_addr_block,
    output[1:0] io_manager_release_bits_payload_client_xact_id,
    output[2:0] io_manager_release_bits_payload_r_type,
    output io_manager_release_bits_payload_voluntary,
    output[127:0] io_manager_release_bits_payload_data
);

  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[1:0] Queue_io_deq_bits_header_src;
  wire[1:0] Queue_io_deq_bits_header_dst;
  wire[25:0] Queue_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_io_deq_bits_payload_client_xact_id;
  wire[1:0] Queue_io_deq_bits_payload_addr_beat;
  wire Queue_io_deq_bits_payload_is_builtin_type;
  wire[2:0] Queue_io_deq_bits_payload_a_type;
  wire[16:0] Queue_io_deq_bits_payload_union;
  wire[127:0] Queue_io_deq_bits_payload_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[1:0] Queue_1_io_deq_bits_header_src;
  wire[1:0] Queue_1_io_deq_bits_header_dst;
  wire[25:0] Queue_1_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_1_io_deq_bits_payload_p_type;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire[1:0] Queue_2_io_deq_bits_header_src;
  wire[1:0] Queue_2_io_deq_bits_header_dst;
  wire[1:0] Queue_2_io_deq_bits_payload_addr_beat;
  wire[25:0] Queue_2_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_2_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_2_io_deq_bits_payload_r_type;
  wire Queue_2_io_deq_bits_payload_voluntary;
  wire[127:0] Queue_2_io_deq_bits_payload_data;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire[1:0] Queue_3_io_deq_bits_header_src;
  wire[1:0] Queue_3_io_deq_bits_header_dst;
  wire[1:0] Queue_3_io_deq_bits_payload_addr_beat;
  wire[1:0] Queue_3_io_deq_bits_payload_client_xact_id;
  wire[3:0] Queue_3_io_deq_bits_payload_manager_xact_id;
  wire Queue_3_io_deq_bits_payload_is_builtin_type;
  wire[3:0] Queue_3_io_deq_bits_payload_g_type;
  wire[127:0] Queue_3_io_deq_bits_payload_data;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_header_src;
  wire[1:0] Queue_4_io_deq_bits_header_dst;
  wire[3:0] Queue_4_io_deq_bits_payload_manager_xact_id;


  assign io_manager_release_bits_payload_data = Queue_2_io_deq_bits_payload_data;
  assign io_manager_release_bits_payload_voluntary = Queue_2_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_2_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_client_xact_id = Queue_2_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_addr_block = Queue_2_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_addr_beat = Queue_2_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_header_dst = Queue_2_io_deq_bits_header_dst;
  assign io_manager_release_bits_header_src = Queue_2_io_deq_bits_header_src;
  assign io_manager_release_valid = Queue_2_io_deq_valid;
  assign io_manager_probe_ready = Queue_1_io_enq_ready;
  assign io_manager_finish_bits_payload_manager_xact_id = Queue_4_io_deq_bits_payload_manager_xact_id;
  assign io_manager_finish_bits_header_dst = Queue_4_io_deq_bits_header_dst;
  assign io_manager_finish_bits_header_src = Queue_4_io_deq_bits_header_src;
  assign io_manager_finish_valid = Queue_4_io_deq_valid;
  assign io_manager_grant_ready = Queue_3_io_enq_ready;
  assign io_manager_acquire_bits_payload_data = Queue_io_deq_bits_payload_data;
  assign io_manager_acquire_bits_payload_union = Queue_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_a_type = Queue_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_block = Queue_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_header_dst = Queue_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_header_src = Queue_io_deq_bits_header_src;
  assign io_manager_acquire_valid = Queue_io_deq_valid;
  assign io_client_release_ready = Queue_2_io_enq_ready;
  assign io_client_probe_bits_payload_p_type = Queue_1_io_deq_bits_payload_p_type;
  assign io_client_probe_bits_payload_addr_block = Queue_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_header_dst = Queue_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_header_src = Queue_1_io_deq_bits_header_src;
  assign io_client_probe_valid = Queue_1_io_deq_valid;
  assign io_client_finish_ready = Queue_4_io_enq_ready;
  assign io_client_grant_bits_payload_data = Queue_3_io_deq_bits_payload_data;
  assign io_client_grant_bits_payload_g_type = Queue_3_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_3_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_3_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_client_xact_id = Queue_3_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_addr_beat = Queue_3_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_header_dst = Queue_3_io_deq_bits_header_dst;
  assign io_client_grant_bits_header_src = Queue_3_io_deq_bits_header_src;
  assign io_client_grant_valid = Queue_3_io_deq_valid;
  assign io_client_acquire_ready = Queue_io_enq_ready;
  Queue_8 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_client_acquire_valid ),
       .io_enq_bits_header_src( io_client_acquire_bits_header_src ),
       .io_enq_bits_header_dst( io_client_acquire_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_client_acquire_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_acquire_bits_payload_client_xact_id ),
       .io_enq_bits_payload_addr_beat( io_client_acquire_bits_payload_addr_beat ),
       .io_enq_bits_payload_is_builtin_type( io_client_acquire_bits_payload_is_builtin_type ),
       .io_enq_bits_payload_a_type( io_client_acquire_bits_payload_a_type ),
       .io_enq_bits_payload_union( io_client_acquire_bits_payload_union ),
       .io_enq_bits_payload_data( io_client_acquire_bits_payload_data ),
       .io_deq_ready( io_manager_acquire_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_header_src( Queue_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_addr_beat( Queue_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_is_builtin_type( Queue_io_deq_bits_payload_is_builtin_type ),
       .io_deq_bits_payload_a_type( Queue_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_union( Queue_io_deq_bits_payload_union ),
       .io_deq_bits_payload_data( Queue_io_deq_bits_payload_data )
       //.io_count(  )
  );
  Queue_9 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( io_manager_probe_valid ),
       .io_enq_bits_header_src( io_manager_probe_bits_header_src ),
       .io_enq_bits_header_dst( io_manager_probe_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_manager_probe_bits_payload_addr_block ),
       .io_enq_bits_payload_p_type( io_manager_probe_bits_payload_p_type ),
       .io_deq_ready( io_client_probe_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_header_src( Queue_1_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_1_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_1_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_p_type( Queue_1_io_deq_bits_payload_p_type )
       //.io_count(  )
  );
  Queue_10 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( io_client_release_valid ),
       .io_enq_bits_header_src( io_client_release_bits_header_src ),
       .io_enq_bits_header_dst( io_client_release_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_client_release_bits_payload_addr_beat ),
       .io_enq_bits_payload_addr_block( io_client_release_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_release_bits_payload_client_xact_id ),
       .io_enq_bits_payload_r_type( io_client_release_bits_payload_r_type ),
       .io_enq_bits_payload_voluntary( io_client_release_bits_payload_voluntary ),
       .io_enq_bits_payload_data( io_client_release_bits_payload_data ),
       .io_deq_ready( io_manager_release_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_header_src( Queue_2_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_2_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_2_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_addr_block( Queue_2_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_2_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_r_type( Queue_2_io_deq_bits_payload_r_type ),
       .io_deq_bits_payload_voluntary( Queue_2_io_deq_bits_payload_voluntary ),
       .io_deq_bits_payload_data( Queue_2_io_deq_bits_payload_data )
       //.io_count(  )
  );
  Queue_11 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( io_manager_grant_valid ),
       .io_enq_bits_header_src( io_manager_grant_bits_header_src ),
       .io_enq_bits_header_dst( io_manager_grant_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_manager_grant_bits_payload_addr_beat ),
       .io_enq_bits_payload_client_xact_id( io_manager_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_manager_xact_id( io_manager_grant_bits_payload_manager_xact_id ),
       .io_enq_bits_payload_is_builtin_type( io_manager_grant_bits_payload_is_builtin_type ),
       .io_enq_bits_payload_g_type( io_manager_grant_bits_payload_g_type ),
       .io_enq_bits_payload_data( io_manager_grant_bits_payload_data ),
       .io_deq_ready( io_client_grant_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_header_src( Queue_3_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_3_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_3_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_client_xact_id( Queue_3_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_manager_xact_id( Queue_3_io_deq_bits_payload_manager_xact_id ),
       .io_deq_bits_payload_is_builtin_type( Queue_3_io_deq_bits_payload_is_builtin_type ),
       .io_deq_bits_payload_g_type( Queue_3_io_deq_bits_payload_g_type ),
       .io_deq_bits_payload_data( Queue_3_io_deq_bits_payload_data )
       //.io_count(  )
  );
  Queue_12 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( io_client_finish_valid ),
       .io_enq_bits_header_src( io_client_finish_bits_header_src ),
       .io_enq_bits_header_dst( io_client_finish_bits_header_dst ),
       .io_enq_bits_payload_manager_xact_id( io_client_finish_bits_payload_manager_xact_id ),
       .io_deq_ready( io_manager_finish_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_manager_xact_id( Queue_4_io_deq_bits_payload_manager_xact_id )
       //.io_count(  )
  );
endmodule

module FinishUnit_1(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [1:0] io_grant_bits_header_src,
    input [1:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [1:0] io_grant_bits_payload_client_xact_id,
    input [3:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input [127:0] io_grant_bits_payload_data,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[1:0] io_refill_bits_client_xact_id,
    output[3:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    output[127:0] io_refill_bits_data,
    input  io_finish_ready,
    output io_finish_valid,
    output[1:0] io_finish_bits_header_src,
    output[1:0] io_finish_bits_header_dst,
    output[3:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[3:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T33;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[3:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[1:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T33 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 2'h1;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = io_grant_valid;
  assign io_grant_ready = T27;
  assign T27 = T28 & io_refill_ready;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_1(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [1:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[1:0] io_client_grant_bits_client_xact_id,
    output[3:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    output[127:0] io_client_grant_bits_data,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_addr_beat,
    input [25:0] io_client_release_bits_addr_block,
    input [1:0] io_client_release_bits_client_xact_id,
    input [2:0] io_client_release_bits_r_type,
    input  io_client_release_bits_voluntary,
    input [127:0] io_client_release_bits_data,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[1:0] io_network_acquire_bits_header_src,
    output[1:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[1:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [1:0] io_network_grant_bits_header_src,
    input [1:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [1:0] io_network_grant_bits_payload_client_xact_id,
    input [3:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[1:0] io_network_finish_bits_header_src,
    output[1:0] io_network_finish_bits_header_dst,
    output[3:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [1:0] io_network_probe_bits_header_src,
    input [1:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[1:0] io_network_release_bits_header_src,
    output[1:0] io_network_release_bits_header_dst,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[1:0] io_network_release_bits_payload_client_xact_id,
    output[2:0] io_network_release_bits_payload_r_type,
    output io_network_release_bits_payload_voluntary,
    output[127:0] io_network_release_bits_payload_data
);

  wire[127:0] rel_with_header_bits_payload_data;
  wire rel_with_header_bits_payload_voluntary;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire[1:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[1:0] rel_with_header_bits_header_dst;
  wire[1:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[1:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[1:0] acq_with_header_bits_header_dst;
  wire[1:0] acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[1:0] finisher_io_refill_bits_client_xact_id;
  wire[3:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_finish_valid;
  wire[1:0] finisher_io_finish_bits_header_src;
  wire[1:0] finisher_io_finish_bits_header_dst;
  wire[3:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 2'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 2'h1;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 2'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 2'h1;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_1 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module FinishUnit_2(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [1:0] io_grant_bits_header_src,
    input [1:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [1:0] io_grant_bits_payload_client_xact_id,
    input [3:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input [127:0] io_grant_bits_payload_data,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[1:0] io_refill_bits_client_xact_id,
    output[3:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    output[127:0] io_refill_bits_data,
    input  io_finish_ready,
    output io_finish_valid,
    output[1:0] io_finish_bits_header_src,
    output[1:0] io_finish_bits_header_dst,
    output[3:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[3:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T33;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[3:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[1:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T33 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 2'h2;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = io_grant_valid;
  assign io_grant_ready = T27;
  assign T27 = T28 & io_refill_ready;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_2(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [1:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[1:0] io_client_grant_bits_client_xact_id,
    output[3:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    output[127:0] io_client_grant_bits_data,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_addr_beat,
    input [25:0] io_client_release_bits_addr_block,
    input [1:0] io_client_release_bits_client_xact_id,
    input [2:0] io_client_release_bits_r_type,
    input  io_client_release_bits_voluntary,
    input [127:0] io_client_release_bits_data,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[1:0] io_network_acquire_bits_header_src,
    output[1:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[1:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [1:0] io_network_grant_bits_header_src,
    input [1:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [1:0] io_network_grant_bits_payload_client_xact_id,
    input [3:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[1:0] io_network_finish_bits_header_src,
    output[1:0] io_network_finish_bits_header_dst,
    output[3:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [1:0] io_network_probe_bits_header_src,
    input [1:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[1:0] io_network_release_bits_header_src,
    output[1:0] io_network_release_bits_header_dst,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[1:0] io_network_release_bits_payload_client_xact_id,
    output[2:0] io_network_release_bits_payload_r_type,
    output io_network_release_bits_payload_voluntary,
    output[127:0] io_network_release_bits_payload_data
);

  wire[127:0] rel_with_header_bits_payload_data;
  wire rel_with_header_bits_payload_voluntary;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire[1:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[1:0] rel_with_header_bits_header_dst;
  wire[1:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[1:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[1:0] acq_with_header_bits_header_dst;
  wire[1:0] acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[1:0] finisher_io_refill_bits_client_xact_id;
  wire[3:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_finish_valid;
  wire[1:0] finisher_io_finish_bits_header_src;
  wire[1:0] finisher_io_finish_bits_header_dst;
  wire[3:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 2'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 2'h2;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 2'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 2'h2;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_2 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module ManagerTileLinkNetworkPort(
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[25:0] io_manager_acquire_bits_addr_block,
    output[1:0] io_manager_acquire_bits_client_xact_id,
    output[1:0] io_manager_acquire_bits_addr_beat,
    output io_manager_acquire_bits_is_builtin_type,
    output[2:0] io_manager_acquire_bits_a_type,
    output[16:0] io_manager_acquire_bits_union,
    output[127:0] io_manager_acquire_bits_data,
    output[1:0] io_manager_acquire_bits_client_id,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_addr_beat,
    input [1:0] io_manager_grant_bits_client_xact_id,
    input [3:0] io_manager_grant_bits_manager_xact_id,
    input  io_manager_grant_bits_is_builtin_type,
    input [3:0] io_manager_grant_bits_g_type,
    input [127:0] io_manager_grant_bits_data,
    input [1:0] io_manager_grant_bits_client_id,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[3:0] io_manager_finish_bits_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [25:0] io_manager_probe_bits_addr_block,
    input [1:0] io_manager_probe_bits_p_type,
    input [1:0] io_manager_probe_bits_client_id,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_addr_beat,
    output[25:0] io_manager_release_bits_addr_block,
    output[1:0] io_manager_release_bits_client_xact_id,
    output[2:0] io_manager_release_bits_r_type,
    output io_manager_release_bits_voluntary,
    output[127:0] io_manager_release_bits_data,
    output[1:0] io_manager_release_bits_client_id,
    output io_network_acquire_ready,
    input  io_network_acquire_valid,
    input [1:0] io_network_acquire_bits_header_src,
    input [1:0] io_network_acquire_bits_header_dst,
    input [25:0] io_network_acquire_bits_payload_addr_block,
    input [1:0] io_network_acquire_bits_payload_client_xact_id,
    input [1:0] io_network_acquire_bits_payload_addr_beat,
    input  io_network_acquire_bits_payload_is_builtin_type,
    input [2:0] io_network_acquire_bits_payload_a_type,
    input [16:0] io_network_acquire_bits_payload_union,
    input [127:0] io_network_acquire_bits_payload_data,
    input  io_network_grant_ready,
    output io_network_grant_valid,
    output[1:0] io_network_grant_bits_header_src,
    output[1:0] io_network_grant_bits_header_dst,
    output[1:0] io_network_grant_bits_payload_addr_beat,
    output[1:0] io_network_grant_bits_payload_client_xact_id,
    output[3:0] io_network_grant_bits_payload_manager_xact_id,
    output io_network_grant_bits_payload_is_builtin_type,
    output[3:0] io_network_grant_bits_payload_g_type,
    output[127:0] io_network_grant_bits_payload_data,
    output io_network_finish_ready,
    input  io_network_finish_valid,
    input [1:0] io_network_finish_bits_header_src,
    input [1:0] io_network_finish_bits_header_dst,
    input [3:0] io_network_finish_bits_payload_manager_xact_id,
    input  io_network_probe_ready,
    output io_network_probe_valid,
    output[1:0] io_network_probe_bits_header_src,
    output[1:0] io_network_probe_bits_header_dst,
    output[25:0] io_network_probe_bits_payload_addr_block,
    output[1:0] io_network_probe_bits_payload_p_type,
    output io_network_release_ready,
    input  io_network_release_valid,
    input [1:0] io_network_release_bits_header_src,
    input [1:0] io_network_release_bits_header_dst,
    input [1:0] io_network_release_bits_payload_addr_beat,
    input [25:0] io_network_release_bits_payload_addr_block,
    input [1:0] io_network_release_bits_payload_client_xact_id,
    input [2:0] io_network_release_bits_payload_r_type,
    input  io_network_release_bits_payload_voluntary,
    input [127:0] io_network_release_bits_payload_data
);

  wire T0;
  wire[1:0] T1;
  wire[25:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  wire[127:0] T7;
  wire[3:0] T8;
  wire T9;
  wire[3:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire T15;
  wire T16;
  wire[127:0] T17;
  wire T18;
  wire[2:0] T19;
  wire[1:0] T20;
  wire[25:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire T26;
  wire T27;
  wire[127:0] T28;
  wire[16:0] T29;
  wire[2:0] T30;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[25:0] T34;
  wire T35;


  assign io_network_release_ready = T0;
  assign T0 = io_manager_release_ready;
  assign io_network_probe_bits_payload_p_type = T1;
  assign T1 = io_manager_probe_bits_p_type;
  assign io_network_probe_bits_payload_addr_block = T2;
  assign T2 = io_manager_probe_bits_addr_block;
  assign io_network_probe_bits_header_dst = T3;
  assign T3 = io_manager_probe_bits_client_id;
  assign io_network_probe_bits_header_src = T4;
  assign T4 = 2'h0;
  assign io_network_probe_valid = T5;
  assign T5 = io_manager_probe_valid;
  assign io_network_finish_ready = T6;
  assign T6 = io_manager_finish_ready;
  assign io_network_grant_bits_payload_data = T7;
  assign T7 = io_manager_grant_bits_data;
  assign io_network_grant_bits_payload_g_type = T8;
  assign T8 = io_manager_grant_bits_g_type;
  assign io_network_grant_bits_payload_is_builtin_type = T9;
  assign T9 = io_manager_grant_bits_is_builtin_type;
  assign io_network_grant_bits_payload_manager_xact_id = T10;
  assign T10 = io_manager_grant_bits_manager_xact_id;
  assign io_network_grant_bits_payload_client_xact_id = T11;
  assign T11 = io_manager_grant_bits_client_xact_id;
  assign io_network_grant_bits_payload_addr_beat = T12;
  assign T12 = io_manager_grant_bits_addr_beat;
  assign io_network_grant_bits_header_dst = T13;
  assign T13 = io_manager_grant_bits_client_id;
  assign io_network_grant_bits_header_src = T14;
  assign T14 = 2'h0;
  assign io_network_grant_valid = T15;
  assign T15 = io_manager_grant_valid;
  assign io_network_acquire_ready = T16;
  assign T16 = io_manager_acquire_ready;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src;
  assign io_manager_release_bits_data = T17;
  assign T17 = io_network_release_bits_payload_data;
  assign io_manager_release_bits_voluntary = T18;
  assign T18 = io_network_release_bits_payload_voluntary;
  assign io_manager_release_bits_r_type = T19;
  assign T19 = io_network_release_bits_payload_r_type;
  assign io_manager_release_bits_client_xact_id = T20;
  assign T20 = io_network_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_addr_block = T21;
  assign T21 = io_network_release_bits_payload_addr_block;
  assign io_manager_release_bits_addr_beat = T22;
  assign T22 = io_network_release_bits_payload_addr_beat;
  assign io_manager_release_valid = T23;
  assign T23 = io_network_release_valid;
  assign io_manager_probe_ready = T24;
  assign T24 = io_network_probe_ready;
  assign io_manager_finish_bits_manager_xact_id = T25;
  assign T25 = io_network_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_valid = T26;
  assign T26 = io_network_finish_valid;
  assign io_manager_grant_ready = T27;
  assign T27 = io_network_grant_ready;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src;
  assign io_manager_acquire_bits_data = T28;
  assign T28 = io_network_acquire_bits_payload_data;
  assign io_manager_acquire_bits_union = T29;
  assign T29 = io_network_acquire_bits_payload_union;
  assign io_manager_acquire_bits_a_type = T30;
  assign T30 = io_network_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_is_builtin_type = T31;
  assign T31 = io_network_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_addr_beat = T32;
  assign T32 = io_network_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_client_xact_id = T33;
  assign T33 = io_network_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_addr_block = T34;
  assign T34 = io_network_acquire_bits_payload_addr_block;
  assign io_manager_acquire_valid = T35;
  assign T35 = io_network_acquire_valid;
endmodule

module Queue_13(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_enq_bits_payload_voluntary,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_r_type,
    output io_deq_bits_payload_voluntary,
    output[127:0] io_deq_bits_payload_data,
    output io_count
);

  wire T23;
  wire[1:0] T0;
  reg  full;
  wire T24;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[127:0] T3;
  wire[165:0] T4;
  reg [165:0] ram [0:0];
  wire[165:0] T5;
  wire[165:0] T6;
  wire[165:0] T7;
  wire[133:0] T8;
  wire[128:0] T9;
  wire[4:0] T10;
  wire[31:0] T11;
  wire[27:0] T12;
  wire[3:0] T13;
  wire T14;
  wire[2:0] T15;
  wire[1:0] T16;
  wire[25:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire empty;
  wire T22;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T23;
  assign T23 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T24 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_data = T3;
  assign T3 = T4[7'h7f:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = {io_enq_bits_payload_voluntary, io_enq_bits_payload_data};
  assign T10 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_r_type};
  assign T11 = {T13, T12};
  assign T12 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_addr_block};
  assign T13 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_voluntary = T14;
  assign T14 = T4[8'h80:8'h80];
  assign io_deq_bits_payload_r_type = T15;
  assign T15 = T4[8'h83:8'h81];
  assign io_deq_bits_payload_client_xact_id = T16;
  assign T16 = T4[8'h85:8'h84];
  assign io_deq_bits_payload_addr_block = T17;
  assign T17 = T4[8'h9f:8'h86];
  assign io_deq_bits_payload_addr_beat = T18;
  assign T18 = T4[8'ha1:8'ha0];
  assign io_deq_bits_header_dst = T19;
  assign T19 = T4[8'ha3:8'ha2];
  assign io_deq_bits_header_src = T20;
  assign T20 = T4[8'ha5:8'ha4];
  assign io_deq_valid = T21;
  assign T21 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module TileLinkEnqueuer_1(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [1:0] io_client_acquire_bits_header_src,
    input [1:0] io_client_acquire_bits_header_dst,
    input [25:0] io_client_acquire_bits_payload_addr_block,
    input [1:0] io_client_acquire_bits_payload_client_xact_id,
    input [1:0] io_client_acquire_bits_payload_addr_beat,
    input  io_client_acquire_bits_payload_is_builtin_type,
    input [2:0] io_client_acquire_bits_payload_a_type,
    input [16:0] io_client_acquire_bits_payload_union,
    input [127:0] io_client_acquire_bits_payload_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_header_src,
    output[1:0] io_client_grant_bits_header_dst,
    output[1:0] io_client_grant_bits_payload_addr_beat,
    output[1:0] io_client_grant_bits_payload_client_xact_id,
    output[3:0] io_client_grant_bits_payload_manager_xact_id,
    output io_client_grant_bits_payload_is_builtin_type,
    output[3:0] io_client_grant_bits_payload_g_type,
    output[127:0] io_client_grant_bits_payload_data,
    output io_client_finish_ready,
    input  io_client_finish_valid,
    input [1:0] io_client_finish_bits_header_src,
    input [1:0] io_client_finish_bits_header_dst,
    input [3:0] io_client_finish_bits_payload_manager_xact_id,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[1:0] io_client_probe_bits_header_src,
    output[1:0] io_client_probe_bits_header_dst,
    output[25:0] io_client_probe_bits_payload_addr_block,
    output[1:0] io_client_probe_bits_payload_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_header_src,
    input [1:0] io_client_release_bits_header_dst,
    input [1:0] io_client_release_bits_payload_addr_beat,
    input [25:0] io_client_release_bits_payload_addr_block,
    input [1:0] io_client_release_bits_payload_client_xact_id,
    input [2:0] io_client_release_bits_payload_r_type,
    input  io_client_release_bits_payload_voluntary,
    input [127:0] io_client_release_bits_payload_data,
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[1:0] io_manager_acquire_bits_header_src,
    output[1:0] io_manager_acquire_bits_header_dst,
    output[25:0] io_manager_acquire_bits_payload_addr_block,
    output[1:0] io_manager_acquire_bits_payload_client_xact_id,
    output[1:0] io_manager_acquire_bits_payload_addr_beat,
    output io_manager_acquire_bits_payload_is_builtin_type,
    output[2:0] io_manager_acquire_bits_payload_a_type,
    output[16:0] io_manager_acquire_bits_payload_union,
    output[127:0] io_manager_acquire_bits_payload_data,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_header_src,
    input [1:0] io_manager_grant_bits_header_dst,
    input [1:0] io_manager_grant_bits_payload_addr_beat,
    input [1:0] io_manager_grant_bits_payload_client_xact_id,
    input [3:0] io_manager_grant_bits_payload_manager_xact_id,
    input  io_manager_grant_bits_payload_is_builtin_type,
    input [3:0] io_manager_grant_bits_payload_g_type,
    input [127:0] io_manager_grant_bits_payload_data,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[1:0] io_manager_finish_bits_header_src,
    output[1:0] io_manager_finish_bits_header_dst,
    output[3:0] io_manager_finish_bits_payload_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [1:0] io_manager_probe_bits_header_src,
    input [1:0] io_manager_probe_bits_header_dst,
    input [25:0] io_manager_probe_bits_payload_addr_block,
    input [1:0] io_manager_probe_bits_payload_p_type,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_header_src,
    output[1:0] io_manager_release_bits_header_dst,
    output[1:0] io_manager_release_bits_payload_addr_beat,
    output[25:0] io_manager_release_bits_payload_addr_block,
    output[1:0] io_manager_release_bits_payload_client_xact_id,
    output[2:0] io_manager_release_bits_payload_r_type,
    output io_manager_release_bits_payload_voluntary,
    output[127:0] io_manager_release_bits_payload_data
);

  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[1:0] Queue_io_deq_bits_header_src;
  wire[1:0] Queue_io_deq_bits_header_dst;
  wire[1:0] Queue_io_deq_bits_payload_addr_beat;
  wire[25:0] Queue_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_io_deq_bits_payload_r_type;
  wire Queue_io_deq_bits_payload_voluntary;
  wire[127:0] Queue_io_deq_bits_payload_data;


  assign io_manager_release_bits_payload_data = Queue_io_deq_bits_payload_data;
  assign io_manager_release_bits_payload_voluntary = Queue_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_client_xact_id = Queue_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_addr_block = Queue_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_addr_beat = Queue_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_header_dst = Queue_io_deq_bits_header_dst;
  assign io_manager_release_bits_header_src = Queue_io_deq_bits_header_src;
  assign io_manager_release_valid = Queue_io_deq_valid;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_client_release_ready = Queue_io_enq_ready;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_acquire_ready = io_manager_acquire_ready;
  Queue_13 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_client_release_valid ),
       .io_enq_bits_header_src( io_client_release_bits_header_src ),
       .io_enq_bits_header_dst( io_client_release_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_client_release_bits_payload_addr_beat ),
       .io_enq_bits_payload_addr_block( io_client_release_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_release_bits_payload_client_xact_id ),
       .io_enq_bits_payload_r_type( io_client_release_bits_payload_r_type ),
       .io_enq_bits_payload_voluntary( io_client_release_bits_payload_voluntary ),
       .io_enq_bits_payload_data( io_client_release_bits_payload_data ),
       .io_deq_ready( io_manager_release_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_header_src( Queue_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_addr_block( Queue_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_r_type( Queue_io_deq_bits_payload_r_type ),
       .io_deq_bits_payload_voluntary( Queue_io_deq_bits_payload_voluntary ),
       .io_deq_bits_payload_data( Queue_io_deq_bits_payload_data )
       //.io_count(  )
  );
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input  io_in_2_bits_payload_is_builtin_type,
    input [2:0] io_in_2_bits_payload_a_type,
    input [16:0] io_in_2_bits_payload_union,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input  io_in_1_bits_payload_is_builtin_type,
    input [2:0] io_in_1_bits_payload_a_type,
    input [16:0] io_in_1_bits_payload_union,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input  io_in_0_bits_payload_is_builtin_type,
    input [2:0] io_in_0_bits_payload_a_type,
    input [16:0] io_in_0_bits_payload_union,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr_block,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[1:0] io_out_bits_payload_addr_beat,
    output io_out_bits_payload_is_builtin_type,
    output[2:0] io_out_bits_payload_a_type,
    output[16:0] io_out_bits_payload_union,
    output[127:0] io_out_bits_payload_data,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T107;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  reg [1:0] lockIdx;
  wire[1:0] T108;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg  locked;
  wire T109;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[1:0] T25;
  reg [1:0] R26;
  wire[1:0] T110;
  wire[1:0] T27;
  wire[127:0] T28;
  wire[127:0] T29;
  wire T30;
  wire[1:0] T31;
  wire T32;
  wire[16:0] T33;
  wire[16:0] T34;
  wire T35;
  wire T36;
  wire[2:0] T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire[25:0] T53;
  wire[25:0] T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R26 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T107 = reset ? 2'h0 : T6;
  assign T6 = T7 ? chosen : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign T108 = reset ? 2'h2 : T10;
  assign T10 = T15 ? T11 : lockIdx;
  assign T11 = T14 ? 2'h0 : T12;
  assign T12 = T13 ? 2'h1 : 2'h2;
  assign T13 = io_in_1_ready & io_in_1_valid;
  assign T14 = io_in_0_ready & io_in_0_valid;
  assign T15 = T17 & T16;
  assign T16 = locked ^ 1'h1;
  assign T17 = T20 & T18;
  assign T18 = io_out_bits_payload_is_builtin_type & T19;
  assign T19 = 3'h3 == io_out_bits_payload_a_type;
  assign T20 = io_out_ready & io_out_valid;
  assign T109 = reset ? 1'h0 : T21;
  assign T21 = T23 ? 1'h0 : T22;
  assign T22 = T15 ? 1'h1 : locked;
  assign T23 = T20 & T24;
  assign T24 = T25 == 2'h0;
  assign T25 = R26 + 2'h1;
  assign T110 = reset ? 2'h0 : T27;
  assign T27 = T17 ? T25 : R26;
  assign io_out_bits_payload_data = T28;
  assign T28 = T32 ? io_in_2_bits_payload_data : T29;
  assign T29 = T30 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T30 = T31[1'h0:1'h0];
  assign T31 = chosen;
  assign T32 = T31[1'h1:1'h1];
  assign io_out_bits_payload_union = T33;
  assign T33 = T36 ? io_in_2_bits_payload_union : T34;
  assign T34 = T35 ? io_in_1_bits_payload_union : io_in_0_bits_payload_union;
  assign T35 = T31[1'h0:1'h0];
  assign T36 = T31[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T37;
  assign T37 = T40 ? io_in_2_bits_payload_a_type : T38;
  assign T38 = T39 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T39 = T31[1'h0:1'h0];
  assign T40 = T31[1'h1:1'h1];
  assign io_out_bits_payload_is_builtin_type = T41;
  assign T41 = T44 ? io_in_2_bits_payload_is_builtin_type : T42;
  assign T42 = T43 ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign T43 = T31[1'h0:1'h0];
  assign T44 = T31[1'h1:1'h1];
  assign io_out_bits_payload_addr_beat = T45;
  assign T45 = T48 ? io_in_2_bits_payload_addr_beat : T46;
  assign T46 = T47 ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign T47 = T31[1'h0:1'h0];
  assign T48 = T31[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T49;
  assign T49 = T52 ? io_in_2_bits_payload_client_xact_id : T50;
  assign T50 = T51 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T51 = T31[1'h0:1'h0];
  assign T52 = T31[1'h1:1'h1];
  assign io_out_bits_payload_addr_block = T53;
  assign T53 = T56 ? io_in_2_bits_payload_addr_block : T54;
  assign T54 = T55 ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign T55 = T31[1'h0:1'h0];
  assign T56 = T31[1'h1:1'h1];
  assign io_out_bits_header_dst = T57;
  assign T57 = T60 ? io_in_2_bits_header_dst : T58;
  assign T58 = T59 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T59 = T31[1'h0:1'h0];
  assign T60 = T31[1'h1:1'h1];
  assign io_out_bits_header_src = T61;
  assign T61 = T64 ? io_in_2_bits_header_src : T62;
  assign T62 = T63 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T63 = T31[1'h0:1'h0];
  assign T64 = T31[1'h1:1'h1];
  assign io_out_valid = T65;
  assign T65 = T68 ? io_in_2_valid : T66;
  assign T66 = T67 ? io_in_1_valid : io_in_0_valid;
  assign T67 = T31[1'h0:1'h0];
  assign T68 = T31[1'h1:1'h1];
  assign io_in_0_ready = T69;
  assign T69 = T70 & io_out_ready;
  assign T70 = locked ? T82 : T71;
  assign T71 = T81 | T72;
  assign T72 = T73 ^ 1'h1;
  assign T73 = T76 | T74;
  assign T74 = io_in_2_valid & T75;
  assign T75 = last_grant < 2'h2;
  assign T76 = T79 | T77;
  assign T77 = io_in_1_valid & T78;
  assign T78 = last_grant < 2'h1;
  assign T79 = io_in_0_valid & T80;
  assign T80 = last_grant < 2'h0;
  assign T81 = last_grant < 2'h0;
  assign T82 = lockIdx == 2'h0;
  assign io_in_1_ready = T83;
  assign T83 = T84 & io_out_ready;
  assign T84 = locked ? T93 : T85;
  assign T85 = T90 | T86;
  assign T86 = T87 ^ 1'h1;
  assign T87 = T88 | io_in_0_valid;
  assign T88 = T89 | T74;
  assign T89 = T79 | T77;
  assign T90 = T92 & T91;
  assign T91 = last_grant < 2'h1;
  assign T92 = T79 ^ 1'h1;
  assign T93 = lockIdx == 2'h1;
  assign io_in_2_ready = T94;
  assign T94 = T95 & io_out_ready;
  assign T95 = locked ? T106 : T96;
  assign T96 = T102 | T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T99 | io_in_1_valid;
  assign T99 = T100 | io_in_0_valid;
  assign T100 = T101 | T74;
  assign T101 = T79 | T77;
  assign T102 = T104 & T103;
  assign T103 = last_grant < 2'h2;
  assign T104 = T105 ^ 1'h1;
  assign T105 = T79 | T77;
  assign T106 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T15) begin
      lockIdx <= T11;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T23) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R26 <= 2'h0;
    end else if(T17) begin
      R26 <= T25;
    end
  end
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_r_type,
    input  io_in_2_bits_payload_voluntary,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_r_type,
    input  io_in_1_bits_payload_voluntary,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_in_0_bits_payload_voluntary,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[1:0] io_out_bits_payload_addr_beat,
    output[25:0] io_out_bits_payload_addr_block,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_r_type,
    output io_out_bits_payload_voluntary,
    output[127:0] io_out_bits_payload_data,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T106;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  reg [1:0] lockIdx;
  wire[1:0] T107;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  reg  locked;
  wire T108;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  reg [1:0] R29;
  wire[1:0] T109;
  wire[1:0] T30;
  wire[127:0] T31;
  wire[127:0] T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[2:0] T40;
  wire[2:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire[25:0] T48;
  wire[25:0] T49;
  wire T50;
  wire T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R29 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T106 = reset ? 2'h0 : T6;
  assign T6 = T7 ? chosen : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign T107 = reset ? 2'h2 : T10;
  assign T10 = T15 ? T11 : lockIdx;
  assign T11 = T14 ? 2'h0 : T12;
  assign T12 = T13 ? 2'h1 : 2'h2;
  assign T13 = io_in_1_ready & io_in_1_valid;
  assign T14 = io_in_0_ready & io_in_0_valid;
  assign T15 = T17 & T16;
  assign T16 = locked ^ 1'h1;
  assign T17 = T23 & T18;
  assign T18 = T20 | T19;
  assign T19 = 3'h2 == io_out_bits_payload_r_type;
  assign T20 = T22 | T21;
  assign T21 = 3'h1 == io_out_bits_payload_r_type;
  assign T22 = 3'h0 == io_out_bits_payload_r_type;
  assign T23 = io_out_ready & io_out_valid;
  assign T108 = reset ? 1'h0 : T24;
  assign T24 = T26 ? 1'h0 : T25;
  assign T25 = T15 ? 1'h1 : locked;
  assign T26 = T23 & T27;
  assign T27 = T28 == 2'h0;
  assign T28 = R29 + 2'h1;
  assign T109 = reset ? 2'h0 : T30;
  assign T30 = T17 ? T28 : R29;
  assign io_out_bits_payload_data = T31;
  assign T31 = T35 ? io_in_2_bits_payload_data : T32;
  assign T32 = T33 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T33 = T34[1'h0:1'h0];
  assign T34 = chosen;
  assign T35 = T34[1'h1:1'h1];
  assign io_out_bits_payload_voluntary = T36;
  assign T36 = T39 ? io_in_2_bits_payload_voluntary : T37;
  assign T37 = T38 ? io_in_1_bits_payload_voluntary : io_in_0_bits_payload_voluntary;
  assign T38 = T34[1'h0:1'h0];
  assign T39 = T34[1'h1:1'h1];
  assign io_out_bits_payload_r_type = T40;
  assign T40 = T43 ? io_in_2_bits_payload_r_type : T41;
  assign T41 = T42 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T42 = T34[1'h0:1'h0];
  assign T43 = T34[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T44;
  assign T44 = T47 ? io_in_2_bits_payload_client_xact_id : T45;
  assign T45 = T46 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T46 = T34[1'h0:1'h0];
  assign T47 = T34[1'h1:1'h1];
  assign io_out_bits_payload_addr_block = T48;
  assign T48 = T51 ? io_in_2_bits_payload_addr_block : T49;
  assign T49 = T50 ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign T50 = T34[1'h0:1'h0];
  assign T51 = T34[1'h1:1'h1];
  assign io_out_bits_payload_addr_beat = T52;
  assign T52 = T55 ? io_in_2_bits_payload_addr_beat : T53;
  assign T53 = T54 ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign T54 = T34[1'h0:1'h0];
  assign T55 = T34[1'h1:1'h1];
  assign io_out_bits_header_dst = T56;
  assign T56 = T59 ? io_in_2_bits_header_dst : T57;
  assign T57 = T58 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T58 = T34[1'h0:1'h0];
  assign T59 = T34[1'h1:1'h1];
  assign io_out_bits_header_src = T60;
  assign T60 = T63 ? io_in_2_bits_header_src : T61;
  assign T61 = T62 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T62 = T34[1'h0:1'h0];
  assign T63 = T34[1'h1:1'h1];
  assign io_out_valid = T64;
  assign T64 = T67 ? io_in_2_valid : T65;
  assign T65 = T66 ? io_in_1_valid : io_in_0_valid;
  assign T66 = T34[1'h0:1'h0];
  assign T67 = T34[1'h1:1'h1];
  assign io_in_0_ready = T68;
  assign T68 = T69 & io_out_ready;
  assign T69 = locked ? T81 : T70;
  assign T70 = T80 | T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T75 | T73;
  assign T73 = io_in_2_valid & T74;
  assign T74 = last_grant < 2'h2;
  assign T75 = T78 | T76;
  assign T76 = io_in_1_valid & T77;
  assign T77 = last_grant < 2'h1;
  assign T78 = io_in_0_valid & T79;
  assign T79 = last_grant < 2'h0;
  assign T80 = last_grant < 2'h0;
  assign T81 = lockIdx == 2'h0;
  assign io_in_1_ready = T82;
  assign T82 = T83 & io_out_ready;
  assign T83 = locked ? T92 : T84;
  assign T84 = T89 | T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T87 | io_in_0_valid;
  assign T87 = T88 | T73;
  assign T88 = T78 | T76;
  assign T89 = T91 & T90;
  assign T90 = last_grant < 2'h1;
  assign T91 = T78 ^ 1'h1;
  assign T92 = lockIdx == 2'h1;
  assign io_in_2_ready = T93;
  assign T93 = T94 & io_out_ready;
  assign T94 = locked ? T105 : T95;
  assign T95 = T101 | T96;
  assign T96 = T97 ^ 1'h1;
  assign T97 = T98 | io_in_1_valid;
  assign T98 = T99 | io_in_0_valid;
  assign T99 = T100 | T73;
  assign T100 = T78 | T76;
  assign T101 = T103 & T102;
  assign T102 = last_grant < 2'h2;
  assign T103 = T104 ^ 1'h1;
  assign T104 = T78 | T76;
  assign T105 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T15) begin
      lockIdx <= T11;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T26) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R29 <= 2'h0;
    end else if(T17) begin
      R29 <= T28;
    end
  end
endmodule

module RRArbiter_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[3:0] io_out_bits_payload_manager_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire T3;
  wire T4;
  reg [1:0] last_grant;
  wire[1:0] T58;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T7 ? 2'h1 : T0;
  assign T0 = T3 ? 2'h2 : T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T3 = io_in_2_valid & T4;
  assign T4 = last_grant < 2'h2;
  assign T58 = reset ? 2'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = io_in_1_valid & T8;
  assign T8 = last_grant < 2'h1;
  assign io_out_bits_payload_manager_xact_id = T9;
  assign T9 = T13 ? io_in_2_bits_payload_manager_xact_id : T10;
  assign T10 = T11 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = chosen;
  assign T13 = T12[1'h1:1'h1];
  assign io_out_bits_header_dst = T14;
  assign T14 = T17 ? io_in_2_bits_header_dst : T15;
  assign T15 = T16 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T16 = T12[1'h0:1'h0];
  assign T17 = T12[1'h1:1'h1];
  assign io_out_bits_header_src = T18;
  assign T18 = T21 ? io_in_2_bits_header_src : T19;
  assign T19 = T20 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign io_out_valid = T22;
  assign T22 = T25 ? io_in_2_valid : T23;
  assign T23 = T24 ? io_in_1_valid : io_in_0_valid;
  assign T24 = T12[1'h0:1'h0];
  assign T25 = T12[1'h1:1'h1];
  assign io_in_0_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T37 | T28;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T32 | T30;
  assign T30 = io_in_2_valid & T31;
  assign T31 = last_grant < 2'h2;
  assign T32 = T35 | T33;
  assign T33 = io_in_1_valid & T34;
  assign T34 = last_grant < 2'h1;
  assign T35 = io_in_0_valid & T36;
  assign T36 = last_grant < 2'h0;
  assign T37 = last_grant < 2'h0;
  assign io_in_1_ready = T38;
  assign T38 = T39 & io_out_ready;
  assign T39 = T44 | T40;
  assign T40 = T41 ^ 1'h1;
  assign T41 = T42 | io_in_0_valid;
  assign T42 = T43 | T30;
  assign T43 = T35 | T33;
  assign T44 = T46 & T45;
  assign T45 = last_grant < 2'h1;
  assign T46 = T35 ^ 1'h1;
  assign io_in_2_ready = T47;
  assign T47 = T48 & io_out_ready;
  assign T48 = T54 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_1_valid;
  assign T51 = T52 | io_in_0_valid;
  assign T52 = T53 | T30;
  assign T53 = T35 | T33;
  assign T54 = T56 & T55;
  assign T55 = last_grant < 2'h2;
  assign T56 = T57 ^ 1'h1;
  assign T57 = T35 | T33;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module RocketChipTileLinkArbiter(input clk, input reset,
    output io_clients_2_acquire_ready,
    input  io_clients_2_acquire_valid,
    input [25:0] io_clients_2_acquire_bits_addr_block,
    input [1:0] io_clients_2_acquire_bits_client_xact_id,
    input [1:0] io_clients_2_acquire_bits_addr_beat,
    input  io_clients_2_acquire_bits_is_builtin_type,
    input [2:0] io_clients_2_acquire_bits_a_type,
    input [16:0] io_clients_2_acquire_bits_union,
    input [127:0] io_clients_2_acquire_bits_data,
    input  io_clients_2_grant_ready,
    output io_clients_2_grant_valid,
    output[1:0] io_clients_2_grant_bits_addr_beat,
    output[1:0] io_clients_2_grant_bits_client_xact_id,
    output[3:0] io_clients_2_grant_bits_manager_xact_id,
    output io_clients_2_grant_bits_is_builtin_type,
    output[3:0] io_clients_2_grant_bits_g_type,
    output[127:0] io_clients_2_grant_bits_data,
    input  io_clients_2_probe_ready,
    output io_clients_2_probe_valid,
    output[25:0] io_clients_2_probe_bits_addr_block,
    output[1:0] io_clients_2_probe_bits_p_type,
    output io_clients_2_release_ready,
    input  io_clients_2_release_valid,
    input [1:0] io_clients_2_release_bits_addr_beat,
    input [25:0] io_clients_2_release_bits_addr_block,
    input [1:0] io_clients_2_release_bits_client_xact_id,
    input [2:0] io_clients_2_release_bits_r_type,
    input  io_clients_2_release_bits_voluntary,
    input [127:0] io_clients_2_release_bits_data,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [25:0] io_clients_1_acquire_bits_addr_block,
    input [1:0] io_clients_1_acquire_bits_client_xact_id,
    input [1:0] io_clients_1_acquire_bits_addr_beat,
    input  io_clients_1_acquire_bits_is_builtin_type,
    input [2:0] io_clients_1_acquire_bits_a_type,
    input [16:0] io_clients_1_acquire_bits_union,
    input [127:0] io_clients_1_acquire_bits_data,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_addr_beat,
    output[1:0] io_clients_1_grant_bits_client_xact_id,
    output[3:0] io_clients_1_grant_bits_manager_xact_id,
    output io_clients_1_grant_bits_is_builtin_type,
    output[3:0] io_clients_1_grant_bits_g_type,
    output[127:0] io_clients_1_grant_bits_data,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[25:0] io_clients_1_probe_bits_addr_block,
    output[1:0] io_clients_1_probe_bits_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [1:0] io_clients_1_release_bits_addr_beat,
    input [25:0] io_clients_1_release_bits_addr_block,
    input [1:0] io_clients_1_release_bits_client_xact_id,
    input [2:0] io_clients_1_release_bits_r_type,
    input  io_clients_1_release_bits_voluntary,
    input [127:0] io_clients_1_release_bits_data,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [25:0] io_clients_0_acquire_bits_addr_block,
    input [1:0] io_clients_0_acquire_bits_client_xact_id,
    input [1:0] io_clients_0_acquire_bits_addr_beat,
    input  io_clients_0_acquire_bits_is_builtin_type,
    input [2:0] io_clients_0_acquire_bits_a_type,
    input [16:0] io_clients_0_acquire_bits_union,
    input [127:0] io_clients_0_acquire_bits_data,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_addr_beat,
    output[1:0] io_clients_0_grant_bits_client_xact_id,
    output[3:0] io_clients_0_grant_bits_manager_xact_id,
    output io_clients_0_grant_bits_is_builtin_type,
    output[3:0] io_clients_0_grant_bits_g_type,
    output[127:0] io_clients_0_grant_bits_data,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[25:0] io_clients_0_probe_bits_addr_block,
    output[1:0] io_clients_0_probe_bits_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [1:0] io_clients_0_release_bits_addr_beat,
    input [25:0] io_clients_0_release_bits_addr_block,
    input [1:0] io_clients_0_release_bits_client_xact_id,
    input [2:0] io_clients_0_release_bits_r_type,
    input  io_clients_0_release_bits_voluntary,
    input [127:0] io_clients_0_release_bits_data,
    input  io_managers_0_acquire_ready,
    output io_managers_0_acquire_valid,
    output[25:0] io_managers_0_acquire_bits_addr_block,
    output[1:0] io_managers_0_acquire_bits_client_xact_id,
    output[1:0] io_managers_0_acquire_bits_addr_beat,
    output io_managers_0_acquire_bits_is_builtin_type,
    output[2:0] io_managers_0_acquire_bits_a_type,
    output[16:0] io_managers_0_acquire_bits_union,
    output[127:0] io_managers_0_acquire_bits_data,
    output[1:0] io_managers_0_acquire_bits_client_id,
    output io_managers_0_grant_ready,
    input  io_managers_0_grant_valid,
    input [1:0] io_managers_0_grant_bits_addr_beat,
    input [1:0] io_managers_0_grant_bits_client_xact_id,
    input [3:0] io_managers_0_grant_bits_manager_xact_id,
    input  io_managers_0_grant_bits_is_builtin_type,
    input [3:0] io_managers_0_grant_bits_g_type,
    input [127:0] io_managers_0_grant_bits_data,
    input [1:0] io_managers_0_grant_bits_client_id,
    input  io_managers_0_finish_ready,
    output io_managers_0_finish_valid,
    output[3:0] io_managers_0_finish_bits_manager_xact_id,
    output io_managers_0_probe_ready,
    input  io_managers_0_probe_valid,
    input [25:0] io_managers_0_probe_bits_addr_block,
    input [1:0] io_managers_0_probe_bits_p_type,
    input [1:0] io_managers_0_probe_bits_client_id,
    input  io_managers_0_release_ready,
    output io_managers_0_release_valid,
    output[1:0] io_managers_0_release_bits_addr_beat,
    output[25:0] io_managers_0_release_bits_addr_block,
    output[1:0] io_managers_0_release_bits_client_xact_id,
    output[2:0] io_managers_0_release_bits_r_type,
    output io_managers_0_release_bits_voluntary,
    output[127:0] io_managers_0_release_bits_data,
    output[1:0] io_managers_0_release_bits_client_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  wire[16:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_manager_grant_ready;
  wire ManagerTileLinkNetworkPort_io_manager_finish_valid;
  wire[3:0] ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_manager_probe_ready;
  wire ManagerTileLinkNetworkPort_io_manager_release_valid;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  wire ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_network_acquire_ready;
  wire ManagerTileLinkNetworkPort_io_network_grant_valid;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_header_src;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id;
  wire[3:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type;
  wire[3:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type;
  wire[127:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data;
  wire ManagerTileLinkNetworkPort_io_network_finish_ready;
  wire ManagerTileLinkNetworkPort_io_network_probe_valid;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_header_src;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst;
  wire[25:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type;
  wire ManagerTileLinkNetworkPort_io_network_release_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[1:0] LockingRRArbiter_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_io_out_bits_payload_addr_block;
  wire[1:0] LockingRRArbiter_io_out_bits_payload_client_xact_id;
  wire[1:0] LockingRRArbiter_io_out_bits_payload_addr_beat;
  wire LockingRRArbiter_io_out_bits_payload_is_builtin_type;
  wire[2:0] LockingRRArbiter_io_out_bits_payload_a_type;
  wire[16:0] LockingRRArbiter_io_out_bits_payload_union;
  wire[127:0] LockingRRArbiter_io_out_bits_payload_data;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_addr_beat;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr_block;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_r_type;
  wire LockingRRArbiter_1_io_out_bits_payload_voluntary;
  wire[127:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire RRArbiter_io_in_2_ready;
  wire RRArbiter_io_in_1_ready;
  wire RRArbiter_io_in_0_ready;
  wire RRArbiter_io_out_valid;
  wire[1:0] RRArbiter_io_out_bits_header_src;
  wire[1:0] RRArbiter_io_out_bits_header_dst;
  wire[3:0] RRArbiter_io_out_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_client_acquire_ready;
  wire TileLinkEnqueuer_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_io_client_finish_ready;
  wire TileLinkEnqueuer_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_io_client_release_ready;
  wire TileLinkEnqueuer_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_io_manager_grant_ready;
  wire TileLinkEnqueuer_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_manager_finish_bits_header_dst;
  wire[3:0] TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_manager_probe_ready;
  wire TileLinkEnqueuer_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_io_manager_release_bits_payload_voluntary;
  wire[127:0] TileLinkEnqueuer_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_1_io_client_acquire_ready;
  wire TileLinkEnqueuer_1_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_1_io_client_finish_ready;
  wire TileLinkEnqueuer_1_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_1_io_client_release_ready;
  wire TileLinkEnqueuer_1_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_1_io_manager_grant_ready;
  wire TileLinkEnqueuer_1_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_1_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_manager_finish_bits_header_dst;
  wire[3:0] TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_manager_probe_ready;
  wire TileLinkEnqueuer_1_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary;
  wire[127:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_2_io_client_acquire_ready;
  wire TileLinkEnqueuer_2_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_2_io_client_finish_ready;
  wire TileLinkEnqueuer_2_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_2_io_client_release_ready;
  wire TileLinkEnqueuer_2_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_2_io_manager_grant_ready;
  wire TileLinkEnqueuer_2_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_2_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_manager_finish_bits_header_dst;
  wire[3:0] TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_2_io_manager_probe_ready;
  wire TileLinkEnqueuer_2_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary;
  wire[127:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_3_io_client_acquire_ready;
  wire TileLinkEnqueuer_3_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_3_io_client_finish_ready;
  wire TileLinkEnqueuer_3_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_3_io_client_release_ready;
  wire TileLinkEnqueuer_3_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_3_io_manager_grant_ready;
  wire TileLinkEnqueuer_3_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_3_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_manager_finish_bits_header_dst;
  wire[3:0] TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_3_io_manager_probe_ready;
  wire TileLinkEnqueuer_3_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary;
  wire[127:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_data;
  wire ClientTileLinkNetworkPort_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  wire[127:0] ClientTileLinkNetworkPort_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_io_client_release_ready;
  wire ClientTileLinkNetworkPort_io_network_acquire_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat;
  wire ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union;
  wire[127:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_io_network_finish_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_network_finish_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_io_network_finish_bits_header_dst;
  wire[3:0] ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_io_network_release_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_header_dst;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat;
  wire[25:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id;
  wire[2:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type;
  wire ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary;
  wire[127:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_data;
  wire ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_1_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire[127:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_1_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_1_io_client_release_ready;
  wire ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire[127:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_1_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_1_io_network_finish_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire[3:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_1_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_1_io_network_release_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire[25:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire[127:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire ClientTileLinkNetworkPort_2_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_2_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type;
  wire[127:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_2_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_2_io_client_release_ready;
  wire ClientTileLinkNetworkPort_2_io_network_acquire_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat;
  wire ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union;
  wire[127:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_2_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_2_io_network_finish_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst;
  wire[3:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_2_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_2_io_network_release_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat;
  wire[25:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type;
  wire ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary;
  wire[127:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data;


  assign T0 = T5 ? TileLinkEnqueuer_2_io_manager_probe_ready : T1;
  assign T1 = T4 ? TileLinkEnqueuer_1_io_manager_probe_ready : T2;
  assign T2 = T3 ? TileLinkEnqueuer_io_manager_probe_ready : 1'h0;
  assign T3 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst == 2'h0;
  assign T4 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst == 2'h1;
  assign T5 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst == 2'h2;
  assign T6 = T11 ? TileLinkEnqueuer_2_io_manager_grant_ready : T7;
  assign T7 = T10 ? TileLinkEnqueuer_1_io_manager_grant_ready : T8;
  assign T8 = T9 ? TileLinkEnqueuer_io_manager_grant_ready : 1'h0;
  assign T9 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst == 2'h0;
  assign T10 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst == 2'h1;
  assign T11 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst == 2'h2;
  assign T12 = T5 ? TileLinkEnqueuer_3_io_client_probe_valid : 1'h0;
  assign T13 = T11 ? TileLinkEnqueuer_3_io_client_grant_valid : 1'h0;
  assign T14 = T4 ? TileLinkEnqueuer_3_io_client_probe_valid : 1'h0;
  assign T15 = T10 ? TileLinkEnqueuer_3_io_client_grant_valid : 1'h0;
  assign T16 = T3 ? TileLinkEnqueuer_3_io_client_probe_valid : 1'h0;
  assign T17 = T9 ? TileLinkEnqueuer_3_io_client_grant_valid : 1'h0;
  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_io_manager_release_valid;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_io_manager_probe_ready;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_io_manager_finish_valid;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_io_manager_grant_ready;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  assign io_clients_0_release_ready = ClientTileLinkNetworkPort_io_client_release_ready;
  assign io_clients_0_probe_bits_p_type = ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  assign io_clients_0_probe_bits_addr_block = ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  assign io_clients_0_probe_valid = ClientTileLinkNetworkPort_io_client_probe_valid;
  assign io_clients_0_grant_bits_data = ClientTileLinkNetworkPort_io_client_grant_bits_data;
  assign io_clients_0_grant_bits_g_type = ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  assign io_clients_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  assign io_clients_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  assign io_clients_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  assign io_clients_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  assign io_clients_0_grant_valid = ClientTileLinkNetworkPort_io_client_grant_valid;
  assign io_clients_0_acquire_ready = ClientTileLinkNetworkPort_io_client_acquire_ready;
  assign io_clients_1_release_ready = ClientTileLinkNetworkPort_1_io_client_release_ready;
  assign io_clients_1_probe_bits_p_type = ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  assign io_clients_1_probe_bits_addr_block = ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  assign io_clients_1_probe_valid = ClientTileLinkNetworkPort_1_io_client_probe_valid;
  assign io_clients_1_grant_bits_data = ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_clients_1_grant_bits_g_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_1_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_1_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_1_grant_bits_client_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_1_grant_bits_addr_beat = ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_1_grant_valid = ClientTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_1_acquire_ready = ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_2_release_ready = ClientTileLinkNetworkPort_2_io_client_release_ready;
  assign io_clients_2_probe_bits_p_type = ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type;
  assign io_clients_2_probe_bits_addr_block = ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block;
  assign io_clients_2_probe_valid = ClientTileLinkNetworkPort_2_io_client_probe_valid;
  assign io_clients_2_grant_bits_data = ClientTileLinkNetworkPort_2_io_client_grant_bits_data;
  assign io_clients_2_grant_bits_g_type = ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type;
  assign io_clients_2_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type;
  assign io_clients_2_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id;
  assign io_clients_2_grant_bits_client_xact_id = ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id;
  assign io_clients_2_grant_bits_addr_beat = ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat;
  assign io_clients_2_grant_valid = ClientTileLinkNetworkPort_2_io_client_grant_valid;
  assign io_clients_2_acquire_ready = ClientTileLinkNetworkPort_2_io_client_acquire_ready;
  ClientTileLinkNetworkPort_0 ClientTileLinkNetworkPort(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_0_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_0_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_0_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_0_acquire_bits_addr_beat ),
       .io_client_acquire_bits_is_builtin_type( io_clients_0_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_0_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_0_acquire_bits_union ),
       .io_client_acquire_bits_data( io_clients_0_acquire_bits_data ),
       .io_client_grant_ready( io_clients_0_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_io_client_grant_bits_g_type ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_io_client_grant_bits_data ),
       .io_client_probe_ready( io_clients_0_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_io_client_release_ready ),
       .io_client_release_valid( io_clients_0_release_valid ),
       .io_client_release_bits_addr_beat( io_clients_0_release_bits_addr_beat ),
       .io_client_release_bits_addr_block( io_clients_0_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_0_release_bits_client_xact_id ),
       .io_client_release_bits_r_type( io_clients_0_release_bits_r_type ),
       .io_client_release_bits_voluntary( io_clients_0_release_bits_voluntary ),
       .io_client_release_bits_data( io_clients_0_release_bits_data ),
       .io_network_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_network_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data )
  );
  TileLinkEnqueuer_0 TileLinkEnqueuer(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data ),
       .io_manager_acquire_ready( LockingRRArbiter_io_in_0_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_io_manager_grant_ready ),
       .io_manager_grant_valid( T17 ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_manager_finish_ready( RRArbiter_io_in_0_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_io_manager_probe_ready ),
       .io_manager_probe_valid( T16 ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_io_manager_release_bits_payload_data )
  );
  ClientTileLinkNetworkPort_1 ClientTileLinkNetworkPort_1(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_1_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_1_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_1_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_1_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_1_acquire_bits_addr_beat ),
       .io_client_acquire_bits_is_builtin_type( io_clients_1_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_1_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_1_acquire_bits_union ),
       .io_client_acquire_bits_data( io_clients_1_acquire_bits_data ),
       .io_client_grant_ready( io_clients_1_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_1_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_1_io_client_grant_bits_data ),
       .io_client_probe_ready( io_clients_1_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_1_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_1_io_client_release_ready ),
       .io_client_release_valid( io_clients_1_release_valid ),
       .io_client_release_bits_addr_beat( io_clients_1_release_bits_addr_beat ),
       .io_client_release_bits_addr_block( io_clients_1_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_1_release_bits_client_xact_id ),
       .io_client_release_bits_r_type( io_clients_1_release_bits_r_type ),
       .io_client_release_bits_voluntary( io_clients_1_release_bits_voluntary ),
       .io_client_release_bits_data( io_clients_1_release_bits_data ),
       .io_network_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_1_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_1_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_network_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_1_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_1_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_1_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_1_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data )
  );
  TileLinkEnqueuer_0 TileLinkEnqueuer_1(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_1_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_1_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_1_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_1_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_1_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_1_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data ),
       .io_manager_acquire_ready( LockingRRArbiter_io_in_1_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_1_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_1_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_1_io_manager_grant_ready ),
       .io_manager_grant_valid( T15 ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_manager_finish_ready( RRArbiter_io_in_1_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_1_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_1_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_1_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_1_io_manager_probe_ready ),
       .io_manager_probe_valid( T14 ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_1_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_1_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_1_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_1_io_manager_release_bits_payload_data )
  );
  ClientTileLinkNetworkPort_2 ClientTileLinkNetworkPort_2(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_2_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_2_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_2_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_2_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_2_acquire_bits_addr_beat ),
       .io_client_acquire_bits_is_builtin_type( io_clients_2_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_2_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_2_acquire_bits_union ),
       .io_client_acquire_bits_data( io_clients_2_acquire_bits_data ),
       .io_client_grant_ready( io_clients_2_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_2_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_2_io_client_grant_bits_data ),
       .io_client_probe_ready( io_clients_2_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_2_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_2_io_client_release_ready ),
       .io_client_release_valid( io_clients_2_release_valid ),
       .io_client_release_bits_addr_beat( io_clients_2_release_bits_addr_beat ),
       .io_client_release_bits_addr_block( io_clients_2_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_2_release_bits_client_xact_id ),
       .io_client_release_bits_r_type( io_clients_2_release_bits_r_type ),
       .io_client_release_bits_voluntary( io_clients_2_release_bits_voluntary ),
       .io_client_release_bits_data( io_clients_2_release_bits_data ),
       .io_network_acquire_ready( TileLinkEnqueuer_2_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_2_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_2_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_2_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_2_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_2_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_2_io_client_grant_bits_payload_data ),
       .io_network_finish_ready( TileLinkEnqueuer_2_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_2_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_2_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_2_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_2_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_2_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_2_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_2_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_2_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data )
  );
  TileLinkEnqueuer_0 TileLinkEnqueuer_2(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_2_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_2_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_2_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_2_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_2_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_2_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_2_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_2_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_2_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_2_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_2_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_2_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_2_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_2_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_2_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_2_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data ),
       .io_manager_acquire_ready( LockingRRArbiter_io_in_2_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_2_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_2_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_2_io_manager_grant_ready ),
       .io_manager_grant_valid( T13 ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_manager_finish_ready( RRArbiter_io_in_2_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_2_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_2_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_2_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_2_io_manager_probe_ready ),
       .io_manager_probe_valid( T12 ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_2_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_2_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_2_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_2_io_manager_release_bits_payload_data )
  );
  ManagerTileLinkNetworkPort ManagerTileLinkNetworkPort(
       .io_manager_acquire_ready( io_managers_0_acquire_ready ),
       .io_manager_acquire_valid( ManagerTileLinkNetworkPort_io_manager_acquire_valid ),
       .io_manager_acquire_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block ),
       .io_manager_acquire_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id ),
       .io_manager_acquire_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat ),
       .io_manager_acquire_bits_is_builtin_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type ),
       .io_manager_acquire_bits_a_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type ),
       .io_manager_acquire_bits_union( ManagerTileLinkNetworkPort_io_manager_acquire_bits_union ),
       .io_manager_acquire_bits_data( ManagerTileLinkNetworkPort_io_manager_acquire_bits_data ),
       .io_manager_acquire_bits_client_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id ),
       .io_manager_grant_ready( ManagerTileLinkNetworkPort_io_manager_grant_ready ),
       .io_manager_grant_valid( io_managers_0_grant_valid ),
       .io_manager_grant_bits_addr_beat( io_managers_0_grant_bits_addr_beat ),
       .io_manager_grant_bits_client_xact_id( io_managers_0_grant_bits_client_xact_id ),
       .io_manager_grant_bits_manager_xact_id( io_managers_0_grant_bits_manager_xact_id ),
       .io_manager_grant_bits_is_builtin_type( io_managers_0_grant_bits_is_builtin_type ),
       .io_manager_grant_bits_g_type( io_managers_0_grant_bits_g_type ),
       .io_manager_grant_bits_data( io_managers_0_grant_bits_data ),
       .io_manager_grant_bits_client_id( io_managers_0_grant_bits_client_id ),
       .io_manager_finish_ready( io_managers_0_finish_ready ),
       .io_manager_finish_valid( ManagerTileLinkNetworkPort_io_manager_finish_valid ),
       .io_manager_finish_bits_manager_xact_id( ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id ),
       .io_manager_probe_ready( ManagerTileLinkNetworkPort_io_manager_probe_ready ),
       .io_manager_probe_valid( io_managers_0_probe_valid ),
       .io_manager_probe_bits_addr_block( io_managers_0_probe_bits_addr_block ),
       .io_manager_probe_bits_p_type( io_managers_0_probe_bits_p_type ),
       .io_manager_probe_bits_client_id( io_managers_0_probe_bits_client_id ),
       .io_manager_release_ready( io_managers_0_release_ready ),
       .io_manager_release_valid( ManagerTileLinkNetworkPort_io_manager_release_valid ),
       .io_manager_release_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat ),
       .io_manager_release_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block ),
       .io_manager_release_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id ),
       .io_manager_release_bits_r_type( ManagerTileLinkNetworkPort_io_manager_release_bits_r_type ),
       .io_manager_release_bits_voluntary( ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary ),
       .io_manager_release_bits_data( ManagerTileLinkNetworkPort_io_manager_release_bits_data ),
       .io_manager_release_bits_client_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_id ),
       .io_network_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_network_acquire_valid( TileLinkEnqueuer_3_io_manager_acquire_valid ),
       .io_network_acquire_bits_header_src( TileLinkEnqueuer_3_io_manager_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data ),
       .io_network_grant_ready( TileLinkEnqueuer_3_io_manager_grant_ready ),
       .io_network_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_network_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_network_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_network_finish_valid( TileLinkEnqueuer_3_io_manager_finish_valid ),
       .io_network_finish_bits_header_src( TileLinkEnqueuer_3_io_manager_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( TileLinkEnqueuer_3_io_manager_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( TileLinkEnqueuer_3_io_manager_probe_ready ),
       .io_network_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_network_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_network_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_network_release_valid( TileLinkEnqueuer_3_io_manager_release_valid ),
       .io_network_release_bits_header_src( TileLinkEnqueuer_3_io_manager_release_bits_header_src ),
       .io_network_release_bits_header_dst( TileLinkEnqueuer_3_io_manager_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_r_type( TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_data( TileLinkEnqueuer_3_io_manager_release_bits_payload_data )
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_3(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_3_io_client_acquire_ready ),
       .io_client_acquire_valid( LockingRRArbiter_io_out_valid ),
       .io_client_acquire_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_client_acquire_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( LockingRRArbiter_io_out_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( LockingRRArbiter_io_out_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( LockingRRArbiter_io_out_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( LockingRRArbiter_io_out_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( LockingRRArbiter_io_out_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( LockingRRArbiter_io_out_bits_payload_union ),
       .io_client_acquire_bits_payload_data( LockingRRArbiter_io_out_bits_payload_data ),
       .io_client_grant_ready( T6 ),
       .io_client_grant_valid( TileLinkEnqueuer_3_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_3_io_client_finish_ready ),
       .io_client_finish_valid( RRArbiter_io_out_valid ),
       .io_client_finish_bits_header_src( RRArbiter_io_out_bits_header_src ),
       .io_client_finish_bits_header_dst( RRArbiter_io_out_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( RRArbiter_io_out_bits_payload_manager_xact_id ),
       .io_client_probe_ready( T0 ),
       .io_client_probe_valid( TileLinkEnqueuer_3_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_3_io_client_release_ready ),
       .io_client_release_valid( LockingRRArbiter_1_io_out_valid ),
       .io_client_release_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_client_release_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( LockingRRArbiter_1_io_out_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( LockingRRArbiter_1_io_out_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( LockingRRArbiter_1_io_out_bits_payload_voluntary ),
       .io_client_release_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_manager_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_3_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_3_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_3_io_manager_grant_ready ),
       .io_manager_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_manager_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_manager_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_3_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_3_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_3_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_3_io_manager_probe_ready ),
       .io_manager_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_manager_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_manager_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_3_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_3_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_3_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_3_io_manager_release_bits_payload_data )
  );
  LockingRRArbiter_0 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( TileLinkEnqueuer_2_io_manager_acquire_valid ),
       .io_in_2_bits_header_src( TileLinkEnqueuer_2_io_manager_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat ),
       .io_in_2_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_a_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_union( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union ),
       .io_in_2_bits_payload_data( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( TileLinkEnqueuer_1_io_manager_acquire_valid ),
       .io_in_1_bits_header_src( TileLinkEnqueuer_1_io_manager_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat ),
       .io_in_1_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_a_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_union( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union ),
       .io_in_1_bits_payload_data( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( TileLinkEnqueuer_io_manager_acquire_valid ),
       .io_in_0_bits_header_src( TileLinkEnqueuer_io_manager_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( TileLinkEnqueuer_io_manager_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat ),
       .io_in_0_bits_payload_is_builtin_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_a_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_union( TileLinkEnqueuer_io_manager_acquire_bits_payload_union ),
       .io_in_0_bits_payload_data( TileLinkEnqueuer_io_manager_acquire_bits_payload_data ),
       .io_out_ready( TileLinkEnqueuer_3_io_client_acquire_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_a_type( LockingRRArbiter_io_out_bits_payload_a_type ),
       .io_out_bits_payload_union( LockingRRArbiter_io_out_bits_payload_union ),
       .io_out_bits_payload_data( LockingRRArbiter_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( TileLinkEnqueuer_2_io_manager_release_valid ),
       .io_in_2_bits_header_src( TileLinkEnqueuer_2_io_manager_release_bits_header_src ),
       .io_in_2_bits_header_dst( TileLinkEnqueuer_2_io_manager_release_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat ),
       .io_in_2_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_r_type( TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type ),
       .io_in_2_bits_payload_voluntary( TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary ),
       .io_in_2_bits_payload_data( TileLinkEnqueuer_2_io_manager_release_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( TileLinkEnqueuer_1_io_manager_release_valid ),
       .io_in_1_bits_header_src( TileLinkEnqueuer_1_io_manager_release_bits_header_src ),
       .io_in_1_bits_header_dst( TileLinkEnqueuer_1_io_manager_release_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat ),
       .io_in_1_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_r_type( TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type ),
       .io_in_1_bits_payload_voluntary( TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary ),
       .io_in_1_bits_payload_data( TileLinkEnqueuer_1_io_manager_release_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( TileLinkEnqueuer_io_manager_release_valid ),
       .io_in_0_bits_header_src( TileLinkEnqueuer_io_manager_release_bits_header_src ),
       .io_in_0_bits_header_dst( TileLinkEnqueuer_io_manager_release_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat ),
       .io_in_0_bits_payload_addr_block( TileLinkEnqueuer_io_manager_release_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_r_type( TileLinkEnqueuer_io_manager_release_bits_payload_r_type ),
       .io_in_0_bits_payload_voluntary( TileLinkEnqueuer_io_manager_release_bits_payload_voluntary ),
       .io_in_0_bits_payload_data( TileLinkEnqueuer_io_manager_release_bits_payload_data ),
       .io_out_ready( TileLinkEnqueuer_3_io_client_release_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_1_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_1_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type ),
       .io_out_bits_payload_voluntary( LockingRRArbiter_1_io_out_bits_payload_voluntary ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  RRArbiter_3 RRArbiter(.clk(clk), .reset(reset),
       .io_in_2_ready( RRArbiter_io_in_2_ready ),
       .io_in_2_valid( TileLinkEnqueuer_2_io_manager_finish_valid ),
       .io_in_2_bits_header_src( TileLinkEnqueuer_2_io_manager_finish_bits_header_src ),
       .io_in_2_bits_header_dst( TileLinkEnqueuer_2_io_manager_finish_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id ),
       .io_in_1_ready( RRArbiter_io_in_1_ready ),
       .io_in_1_valid( TileLinkEnqueuer_1_io_manager_finish_valid ),
       .io_in_1_bits_header_src( TileLinkEnqueuer_1_io_manager_finish_bits_header_src ),
       .io_in_1_bits_header_dst( TileLinkEnqueuer_1_io_manager_finish_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id ),
       .io_in_0_ready( RRArbiter_io_in_0_ready ),
       .io_in_0_valid( TileLinkEnqueuer_io_manager_finish_valid ),
       .io_in_0_bits_header_src( TileLinkEnqueuer_io_manager_finish_bits_header_src ),
       .io_in_0_bits_header_dst( TileLinkEnqueuer_io_manager_finish_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id ),
       .io_out_ready( TileLinkEnqueuer_3_io_client_finish_ready ),
       .io_out_valid( RRArbiter_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( RRArbiter_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
endmodule

module BroadcastVoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[25:0] io_inner_probe_bits_addr_block
    //output[1:0] io_inner_probe_bits_p_type
    //output[1:0] io_inner_probe_bits_client_id
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [1:0] state;
  wire[1:0] T133;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire oacq_data_done;
  wire T15;
  wire T16;
  wire T17;
  reg [1:0] R18;
  wire[1:0] T134;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire[3:0] T35;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire[1:0] T41;
  wire T42;
  reg  collect_irel_data;
  wire T135;
  wire T43;
  wire T44;
  wire T45;
  wire irel_data_done;
  wire T46;
  wire T47;
  wire T48;
  reg [1:0] R49;
  wire[1:0] T136;
  wire[1:0] T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire[3:0] T65;
  wire[1:0] T66;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T67;
  wire[3:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[1:0] T74;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T75;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T76;
  wire[3:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T82;
  wire[3:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire[16:0] T90;
  wire[16:0] T91;
  wire[15:0] T92;
  wire[2:0] T93;
  wire T94;
  wire[1:0] T95;
  wire[3:0] T137;
  wire[1:0] T96;
  wire[25:0] T97;
  reg [25:0] xact_addr_block;
  wire[25:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  reg [3:0] irel_data_valid;
  wire[3:0] T138;
  wire[3:0] T107;
  wire[3:0] T108;
  wire[3:0] T109;
  wire[3:0] T110;
  wire[3:0] T111;
  wire[3:0] T139;
  wire T112;
  wire[3:0] T113;
  wire[3:0] T114;
  wire[3:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[1:0] T123;
  reg [1:0] xact_client_id;
  wire[1:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire T127;
  wire[3:0] T128;
  wire[1:0] T129;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    R18 = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    collect_irel_data = {1{$random}};
    R49 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_addr_block = {1{$random}};
    irel_data_valid = {1{$random}};
    xact_client_id = {1{$random}};
    xact_client_xact_id = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_inner_probe_bits_client_id = {1{$random}};
//  assign io_inner_probe_bits_p_type = {1{$random}};
//  assign io_inner_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign io_has_release_match = io_inner_release_bits_voluntary;
  assign io_has_acquire_match = 1'h0;
  assign io_has_acquire_conflict = 1'h0;
  assign io_outer_grant_ready = T0;
  assign T0 = T1 ? io_inner_grant_ready : 1'h0;
  assign T1 = 2'h2 == state;
  assign T133 = reset ? 2'h0 : T2;
  assign T2 = T31 ? 2'h0 : T3;
  assign T3 = T29 ? T25 : T4;
  assign T4 = T14 ? 2'h2 : T5;
  assign T5 = T12 ? T6 : state;
  assign T6 = T7 ? 2'h1 : 2'h3;
  assign T7 = T9 | T8;
  assign T8 = 3'h2 == io_inner_release_bits_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h1 == io_inner_release_bits_r_type;
  assign T11 = 3'h0 == io_inner_release_bits_r_type;
  assign T12 = T13 & io_inner_release_valid;
  assign T13 = 2'h0 == state;
  assign T14 = T24 & oacq_data_done;
  assign oacq_data_done = T22 ? T16 : T15;
  assign T15 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T16 = T21 & T17;
  assign T17 = R18 == 2'h3;
  assign T134 = reset ? 2'h0 : T19;
  assign T19 = T21 ? T20 : R18;
  assign T20 = R18 + 2'h1;
  assign T21 = T15 & T22;
  assign T22 = io_outer_acquire_bits_is_builtin_type & T23;
  assign T23 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T24 = 2'h1 == state;
  assign T25 = T26 ? 2'h3 : 2'h0;
  assign T26 = T27 ^ 1'h1;
  assign T27 = io_inner_grant_bits_is_builtin_type & T28;
  assign T28 = io_inner_grant_bits_g_type == 4'h0;
  assign T29 = T1 & T30;
  assign T30 = io_inner_grant_ready & io_inner_grant_valid;
  assign T31 = T32 & io_inner_finish_valid;
  assign T32 = 2'h3 == state;
  assign io_outer_acquire_bits_data = T33;
  assign T33 = T34;
  assign T34 = T89 ? T75 : T35;
  assign T35 = T73 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T36 = T63 ? io_inner_release_bits_data : T37;
  assign T37 = T38 ? io_inner_release_bits_data : xact_data_buffer_0;
  assign T38 = T42 & T39;
  assign T39 = T40[1'h0:1'h0];
  assign T40 = 1'h1 << T41;
  assign T41 = io_inner_release_bits_addr_beat;
  assign T42 = collect_irel_data & io_inner_release_valid;
  assign T135 = reset ? 1'h0 : T43;
  assign T43 = T12 ? T58 : T44;
  assign T44 = T45 ? 1'h0 : collect_irel_data;
  assign T45 = collect_irel_data & irel_data_done;
  assign irel_data_done = T53 ? T47 : T46;
  assign T46 = io_inner_release_ready & io_inner_release_valid;
  assign T47 = T52 & T48;
  assign T48 = R49 == 2'h3;
  assign T136 = reset ? 2'h0 : T50;
  assign T50 = T52 ? T51 : R49;
  assign T51 = R49 + 2'h1;
  assign T52 = T46 & T53;
  assign T53 = T55 | T54;
  assign T54 = 3'h2 == io_inner_release_bits_r_type;
  assign T55 = T57 | T56;
  assign T56 = 3'h1 == io_inner_release_bits_r_type;
  assign T57 = 3'h0 == io_inner_release_bits_r_type;
  assign T58 = T60 | T59;
  assign T59 = 3'h2 == io_inner_release_bits_r_type;
  assign T60 = T62 | T61;
  assign T61 = 3'h1 == io_inner_release_bits_r_type;
  assign T62 = 3'h0 == io_inner_release_bits_r_type;
  assign T63 = T12 & T64;
  assign T64 = T65[1'h0:1'h0];
  assign T65 = 1'h1 << T66;
  assign T66 = 2'h0;
  assign T67 = T71 ? io_inner_release_bits_data : T68;
  assign T68 = T69 ? io_inner_release_bits_data : xact_data_buffer_1;
  assign T69 = T42 & T70;
  assign T70 = T40[1'h1:1'h1];
  assign T71 = T12 & T72;
  assign T72 = T65[1'h1:1'h1];
  assign T73 = T74[1'h0:1'h0];
  assign T74 = oacq_data_cnt;
  assign oacq_data_cnt = T22 ? R18 : 2'h0;
  assign T75 = T88 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T76 = T80 ? io_inner_release_bits_data : T77;
  assign T77 = T78 ? io_inner_release_bits_data : xact_data_buffer_2;
  assign T78 = T42 & T79;
  assign T79 = T40[2'h2:2'h2];
  assign T80 = T12 & T81;
  assign T81 = T65[2'h2:2'h2];
  assign T82 = T86 ? io_inner_release_bits_data : T83;
  assign T83 = T84 ? io_inner_release_bits_data : xact_data_buffer_3;
  assign T84 = T42 & T85;
  assign T85 = T40[2'h3:2'h3];
  assign T86 = T12 & T87;
  assign T87 = T65[2'h3:2'h3];
  assign T88 = T74[1'h0:1'h0];
  assign T89 = T74[1'h1:1'h1];
  assign io_outer_acquire_bits_union = T90;
  assign T90 = T91;
  assign T91 = {T92, 1'h1};
  assign T92 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T93;
  assign T93 = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T94;
  assign T94 = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T95;
  assign T95 = oacq_data_cnt;
  assign io_outer_acquire_bits_client_xact_id = T137;
  assign T137 = {2'h0, T96};
  assign T96 = 2'h0;
  assign io_outer_acquire_bits_addr_block = T97;
  assign T97 = xact_addr_block;
  assign T98 = T12 ? io_inner_release_bits_addr_block : xact_addr_block;
  assign io_outer_acquire_valid = T99;
  assign T99 = T24 ? T100 : 1'h0;
  assign T100 = T121 | T101;
  assign T101 = T106 & T102;
  assign T102 = T103 - 1'h1;
  assign T103 = 1'h1 << T104;
  assign T104 = T105 + 2'h1;
  assign T105 = oacq_data_cnt - oacq_data_cnt;
  assign T106 = irel_data_valid >> oacq_data_cnt;
  assign T138 = reset ? 4'h0 : T107;
  assign T107 = T12 ? T115 : T108;
  assign T108 = T42 ? T109 : irel_data_valid;
  assign T109 = T113 | T110;
  assign T110 = T139 & T111;
  assign T111 = 1'h1 << io_inner_release_bits_addr_beat;
  assign T139 = T112 ? 4'hf : 4'h0;
  assign T112 = 1'h1;
  assign T113 = irel_data_valid & T114;
  assign T114 = ~ T111;
  assign T115 = T116 << io_inner_release_bits_addr_beat;
  assign T116 = T118 | T117;
  assign T117 = 3'h2 == io_inner_release_bits_r_type;
  assign T118 = T120 | T119;
  assign T119 = 3'h1 == io_inner_release_bits_r_type;
  assign T120 = 3'h0 == io_inner_release_bits_r_type;
  assign T121 = collect_irel_data ^ 1'h1;
  assign io_inner_release_ready = T122;
  assign T122 = T13 ? 1'h1 : collect_irel_data;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_finish_ready = T32;
  assign io_inner_grant_bits_client_id = T123;
  assign T123 = xact_client_id;
  assign T124 = T12 ? io_inner_release_bits_client_id : xact_client_id;
  assign io_inner_grant_bits_data = T125;
  assign T125 = 4'h0;
  assign io_inner_grant_bits_g_type = T126;
  assign T126 = 4'h0;
  assign io_inner_grant_bits_is_builtin_type = T127;
  assign T127 = 1'h1;
  assign io_inner_grant_bits_manager_xact_id = T128;
  assign T128 = 4'h0;
  assign io_inner_grant_bits_client_xact_id = T129;
  assign T129 = xact_client_xact_id;
  assign T130 = T12 ? io_inner_release_bits_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T131;
  assign T131 = 2'h0;
  assign io_inner_grant_valid = T132;
  assign T132 = T1 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T31) begin
      state <= 2'h0;
    end else if(T29) begin
      state <= T25;
    end else if(T14) begin
      state <= 2'h2;
    end else if(T12) begin
      state <= T6;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T21) begin
      R18 <= T20;
    end
    if(T63) begin
      xact_data_buffer_0 <= io_inner_release_bits_data;
    end else if(T38) begin
      xact_data_buffer_0 <= io_inner_release_bits_data;
    end
    if(reset) begin
      collect_irel_data <= 1'h0;
    end else if(T12) begin
      collect_irel_data <= T58;
    end else if(T45) begin
      collect_irel_data <= 1'h0;
    end
    if(reset) begin
      R49 <= 2'h0;
    end else if(T52) begin
      R49 <= T51;
    end
    if(T71) begin
      xact_data_buffer_1 <= io_inner_release_bits_data;
    end else if(T69) begin
      xact_data_buffer_1 <= io_inner_release_bits_data;
    end
    if(T80) begin
      xact_data_buffer_2 <= io_inner_release_bits_data;
    end else if(T78) begin
      xact_data_buffer_2 <= io_inner_release_bits_data;
    end
    if(T86) begin
      xact_data_buffer_3 <= io_inner_release_bits_data;
    end else if(T84) begin
      xact_data_buffer_3 <= io_inner_release_bits_data;
    end
    if(T12) begin
      xact_addr_block <= io_inner_release_bits_addr_block;
    end
    if(reset) begin
      irel_data_valid <= 4'h0;
    end else if(T12) begin
      irel_data_valid <= T115;
    end else if(T42) begin
      irel_data_valid <= T109;
    end
    if(T12) begin
      xact_client_id <= io_inner_release_bits_client_id;
    end
    if(T12) begin
      xact_client_xact_id <= io_inner_release_bits_client_xact_id;
    end
  end
endmodule

module BroadcastAcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T400;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T401;
  wire[2:0] T25;
  wire[2:0] T402;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire pending_outer_write_;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[3:0] mask_incoherent;
  wire[3:0] T403;
  wire T51;
  wire T52;
  wire[3:0] mask_self;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T404;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T405;
  wire T58;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[2:0] T62;
  wire pending_outer_read;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire pending_outer_write;
  wire T69;
  wire T70;
  reg [2:0] xact_a_type;
  wire[2:0] T71;
  wire T72;
  wire T73;
  wire T74;
  reg  xact_is_builtin_type;
  wire T75;
  wire T76;
  wire T77;
  reg  release_count;
  wire T406;
  wire[2:0] T407;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T408;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire T85;
  wire[1:0] T409;
  wire T86;
  wire[2:0] T410;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T411;
  wire T90;
  wire T91;
  wire[2:0] T412;
  wire T92;
  wire[2:0] T413;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire oacq_data_done;
  wire T104;
  wire T105;
  wire T106;
  reg [1:0] R107;
  wire[1:0] T414;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire[2:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire ignt_data_done;
  wire T130;
  wire T131;
  wire T132;
  reg [1:0] R133;
  wire[1:0] T415;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire[2:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  reg[0:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire T159;
  reg  collect_iacq_data;
  wire T416;
  wire T160;
  wire T161;
  wire T162;
  wire iacq_data_done;
  wire T163;
  wire T164;
  wire T165;
  reg [1:0] R166;
  wire[1:0] T417;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  reg[0:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  reg [1:0] xact_client_id;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  reg[0:0] T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  reg [25:0] xact_addr_block;
  wire[25:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  reg  pending_ognt_ack;
  wire T418;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[3:0] T214;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[3:0] T220;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T221;
  wire[3:0] T222;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T223;
  wire[3:0] T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[1:0] T228;
  wire T229;
  wire T230;
  wire T231;
  wire[3:0] T232;
  wire[1:0] T233;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T234;
  wire[3:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[1:0] T241;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T242;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T243;
  wire[3:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T249;
  wire[3:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] oacq_write_beat_data;
  wire T257;
  wire[3:0] oacq_probe_data;
  wire T258;
  wire[16:0] T259;
  wire[16:0] T260;
  wire[16:0] T261;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T419;
  wire[12:0] T262;
  wire[6:0] T263;
  wire[2:0] T264;
  reg [16:0] xact_union;
  wire[16:0] T265;
  wire[3:0] T266;
  wire[16:0] T267;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T268;
  wire[15:0] T269;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T270;
  wire[15:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[15:0] T279;
  wire[15:0] T280;
  wire[7:0] T281;
  wire[7:0] T420;
  wire T282;
  wire[1:0] T283;
  wire T284;
  wire[3:0] T285;
  wire[7:0] T286;
  wire[7:0] T421;
  wire T287;
  wire T288;
  wire T289;
  wire[16:0] oacq_probe_union;
  wire[16:0] T290;
  wire[15:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[2:0] T294;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T295;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T296;
  wire T297;
  wire T298;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T299;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T303;
  wire[1:0] T304;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T308;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T309;
  wire[25:0] T310;
  wire[25:0] T311;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T312;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire[1:0] T321;
  wire T322;
  reg [3:0] iacq_data_valid;
  wire[3:0] T422;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[3:0] T326;
  wire[3:0] T327;
  wire[3:0] T423;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire[1:0] T349;
  wire[1:0] T424;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[1:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[25:0] T372;
  wire T373;
  wire T374;
  reg  pending_probes;
  wire T425;
  wire[3:0] T426;
  wire[3:0] T350;
  wire[3:0] T351;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[1:0] T352;
  wire T353;
  wire T354;
  wire[1:0] T429;
  wire T355;
  wire[1:0] T375;
  wire[3:0] T376;
  wire[3:0] T377;
  wire[3:0] T430;
  wire[2:0] T378;
  wire[2:0] T431;
  wire[1:0] T379;
  wire T380;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] T384;
  wire[2:0] T385;
  wire[2:0] T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[3:0] T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire T397;
  wire T398;
  wire T399;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R107 = {1{$random}};
    R133 = {1{$random}};
    T151 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R166 = {1{$random}};
    T175 = 1'b0;
    xact_client_id = {1{$random}};
    T185 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T400 = reset ? 3'h0 : T11;
  assign T11 = T149 ? 3'h0 : T12;
  assign T12 = T147 ? T143 : T13;
  assign T13 = T129 ? T125 : T14;
  assign T14 = T122 ? 3'h5 : T15;
  assign T15 = T120 ? T119 : T16;
  assign T16 = T117 ? T115 : T17;
  assign T17 = T76 ? T61 : T18;
  assign T18 = T59 ? T19 : state;
  assign T19 = T50 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T44 ? T41 : T22;
  assign T22 = T40 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T401;
  assign T401 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T402;
  assign T402 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T39 ? 3'h4 : T29;
  assign T29 = T38 ? 3'h5 : T30;
  assign T30 = T37 ? 3'h3 : T31;
  assign T31 = T36 ? 3'h3 : T32;
  assign T32 = T35 ? 3'h4 : T33;
  assign T33 = T34 ? 3'h1 : 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h5;
  assign T35 = io_inner_acquire_bits_a_type == 3'h4;
  assign T36 = io_inner_acquire_bits_a_type == 3'h3;
  assign T37 = io_inner_acquire_bits_a_type == 3'h2;
  assign T38 = io_inner_acquire_bits_a_type == 3'h1;
  assign T39 = io_inner_acquire_bits_a_type == 3'h0;
  assign T40 = 4'h0 == T24;
  assign T41 = T43 | T42;
  assign T42 = 4'h4 == T24;
  assign T43 = 4'h5 == T24;
  assign T44 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T45;
  assign T45 = T47 | T46;
  assign T46 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T49 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T50 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T403;
  assign T403 = {3'h0, T51};
  assign T51 = ~ T52;
  assign T52 = io_incoherent_0;
  assign mask_self = T56 | T53;
  assign T53 = T404 & T54;
  assign T54 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T404 = T55 ? 4'hf : 4'h0;
  assign T55 = 1'h0;
  assign T56 = T405 & T57;
  assign T57 = ~ T54;
  assign T405 = {3'h0, T58};
  assign T58 = 1'h1;
  assign T59 = T60 & io_inner_acquire_valid;
  assign T60 = 3'h0 == state;
  assign T61 = pending_outer_write ? 3'h3 : T62;
  assign T62 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T66 : T63;
  assign T63 = T65 | T64;
  assign T64 = 4'h1 == io_inner_grant_bits_g_type;
  assign T65 = 4'h0 == io_inner_grant_bits_g_type;
  assign T66 = T68 | T67;
  assign T67 = 4'h4 == io_inner_grant_bits_g_type;
  assign T68 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T69;
  assign T69 = T72 | T70;
  assign T70 = 3'h4 == xact_a_type;
  assign T71 = T59 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T72 = T74 | T73;
  assign T73 = 3'h3 == xact_a_type;
  assign T74 = 3'h2 == xact_a_type;
  assign T75 = T59 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T76 = T103 & T77;
  assign T77 = release_count == 1'h1;
  assign T406 = T407[1'h0:1'h0];
  assign T407 = reset ? 3'h0 : T78;
  assign T78 = T94 ? T413 : T79;
  assign T79 = T103 ? T412 : T80;
  assign T80 = T91 ? T81 : T408;
  assign T408 = {2'h0, release_count};
  assign T81 = T410 + T82;
  assign T82 = {1'h0, T83};
  assign T83 = T409 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = mask_incoherent[2'h3:2'h3];
  assign T409 = {1'h0, T86};
  assign T86 = mask_incoherent[2'h2:2'h2];
  assign T410 = {1'h0, T87};
  assign T87 = T411 + T88;
  assign T88 = {1'h0, T89};
  assign T89 = mask_incoherent[1'h1:1'h1];
  assign T411 = {1'h0, T90};
  assign T90 = mask_incoherent[1'h0:1'h0];
  assign T91 = T59 & T50;
  assign T412 = {2'h0, T92};
  assign T92 = release_count - 1'h1;
  assign T413 = {2'h0, T93};
  assign T93 = release_count - 1'h1;
  assign T94 = T101 & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = T98 | T97;
  assign T97 = 3'h2 == io_inner_release_bits_r_type;
  assign T98 = T100 | T99;
  assign T99 = 3'h1 == io_inner_release_bits_r_type;
  assign T100 = 3'h0 == io_inner_release_bits_r_type;
  assign T101 = T102 & io_inner_release_valid;
  assign T102 = 3'h1 == state;
  assign T103 = T113 & oacq_data_done;
  assign oacq_data_done = T111 ? T105 : T104;
  assign T104 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T105 = T110 & T106;
  assign T106 = R107 == 2'h3;
  assign T414 = reset ? 2'h0 : T108;
  assign T108 = T110 ? T109 : R107;
  assign T109 = R107 + 2'h1;
  assign T110 = T104 & T111;
  assign T111 = io_outer_acquire_bits_is_builtin_type & T112;
  assign T112 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T113 = T114 & io_outer_acquire_ready;
  assign T114 = T101 & T96;
  assign T115 = pending_outer_write ? 3'h3 : T116;
  assign T116 = pending_outer_read ? 3'h2 : 3'h4;
  assign T117 = T94 & T118;
  assign T118 = release_count == 1'h1;
  assign T119 = pending_outer_read ? 3'h2 : 3'h5;
  assign T120 = T121 & oacq_data_done;
  assign T121 = 3'h3 == state;
  assign T122 = T124 & T123;
  assign T123 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T124 = 3'h2 == state;
  assign T125 = T126 ? 3'h6 : 3'h0;
  assign T126 = T127 ^ 1'h1;
  assign T127 = io_inner_grant_bits_is_builtin_type & T128;
  assign T128 = io_inner_grant_bits_g_type == 4'h0;
  assign T129 = T142 & ignt_data_done;
  assign ignt_data_done = T137 ? T131 : T130;
  assign T130 = io_inner_grant_ready & io_inner_grant_valid;
  assign T131 = T136 & T132;
  assign T132 = R133 == 2'h3;
  assign T415 = reset ? 2'h0 : T134;
  assign T134 = T136 ? T135 : R133;
  assign T135 = R133 + 2'h1;
  assign T136 = T130 & T137;
  assign T137 = io_inner_grant_bits_is_builtin_type ? T141 : T138;
  assign T138 = T140 | T139;
  assign T139 = 4'h1 == io_inner_grant_bits_g_type;
  assign T140 = 4'h0 == io_inner_grant_bits_g_type;
  assign T141 = 4'h5 == io_inner_grant_bits_g_type;
  assign T142 = 3'h5 == state;
  assign T143 = T144 ? 3'h6 : 3'h0;
  assign T144 = T145 ^ 1'h1;
  assign T145 = io_inner_grant_bits_is_builtin_type & T146;
  assign T146 = io_inner_grant_bits_g_type == 4'h0;
  assign T147 = T148 & io_inner_grant_ready;
  assign T148 = 3'h4 == state;
  assign T149 = T150 & io_inner_finish_valid;
  assign T150 = 3'h6 == state;
  assign T152 = T153 | reset;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T157 & T155;
  assign T155 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T156 = T59 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T157 = T159 & T158;
  assign T158 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T159 = T174 & collect_iacq_data;
  assign T416 = reset ? 1'h0 : T160;
  assign T160 = T59 ? T172 : T161;
  assign T161 = T162 ? 1'h0 : collect_iacq_data;
  assign T162 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T170 ? T164 : T163;
  assign T163 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T164 = T169 & T165;
  assign T165 = R166 == 2'h3;
  assign T417 = reset ? 2'h0 : T167;
  assign T167 = T169 ? T168 : R166;
  assign T168 = R166 + 2'h1;
  assign T169 = T163 & T170;
  assign T170 = io_inner_acquire_bits_is_builtin_type & T171;
  assign T171 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = state != 3'h0;
  assign T176 = T177 | reset;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T181 & T179;
  assign T179 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T180 = T59 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T181 = T183 & T182;
  assign T182 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T183 = T184 & collect_iacq_data;
  assign T184 = state != 3'h0;
  assign T186 = T187 | reset;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T192 & T189;
  assign T189 = T191 | T190;
  assign T190 = 3'h5 == xact_a_type;
  assign T191 = 3'h4 == xact_a_type;
  assign T192 = T193 & xact_is_builtin_type;
  assign T193 = state != 3'h0;
  assign io_has_release_match = T194;
  assign T194 = T196 & T195;
  assign T195 = state == 3'h1;
  assign T196 = T198 & T197;
  assign T197 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T198 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T199 = T59 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T200;
  assign T200 = T201 & collect_iacq_data;
  assign T201 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T202;
  assign T202 = T204 & T203;
  assign T203 = collect_iacq_data ^ 1'h1;
  assign T204 = T206 & T205;
  assign T205 = state != 3'h0;
  assign T206 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T207;
  assign T207 = T142 ? io_inner_grant_ready : pending_ognt_ack;
  assign T418 = reset ? 1'h0 : T208;
  assign T208 = T120 ? 1'h1 : T209;
  assign T209 = T103 ? 1'h1 : T210;
  assign T210 = T211 ? 1'h0 : pending_ognt_ack;
  assign T211 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T212;
  assign T212 = T258 ? oacq_probe_data : T213;
  assign T213 = T257 ? T220 : T214;
  assign T214 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T215;
  assign T215 = T217 | T216;
  assign T216 = 3'h4 == xact_a_type;
  assign T217 = T219 | T218;
  assign T218 = 3'h0 == xact_a_type;
  assign T219 = 3'h2 == xact_a_type;
  assign T220 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T221;
  assign T221 = T256 ? T242 : T222;
  assign T222 = T240 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T223 = T230 ? io_inner_acquire_bits_data : T224;
  assign T224 = T225 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T225 = T229 & T226;
  assign T226 = T227[1'h0:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = io_inner_acquire_bits_addr_beat;
  assign T229 = collect_iacq_data & io_inner_acquire_valid;
  assign T230 = T59 & T231;
  assign T231 = T232[1'h0:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = 2'h0;
  assign T234 = T238 ? io_inner_acquire_bits_data : T235;
  assign T235 = T236 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T236 = T229 & T237;
  assign T237 = T227[1'h1:1'h1];
  assign T238 = T59 & T239;
  assign T239 = T232[1'h1:1'h1];
  assign T240 = T241[1'h0:1'h0];
  assign T241 = oacq_data_cnt;
  assign oacq_data_cnt = T111 ? R107 : 2'h0;
  assign T242 = T255 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T243 = T247 ? io_inner_acquire_bits_data : T244;
  assign T244 = T245 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T245 = T229 & T246;
  assign T246 = T227[2'h2:2'h2];
  assign T247 = T59 & T248;
  assign T248 = T232[2'h2:2'h2];
  assign T249 = T253 ? io_inner_acquire_bits_data : T250;
  assign T250 = T251 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T251 = T229 & T252;
  assign T252 = T227[2'h3:2'h3];
  assign T253 = T59 & T254;
  assign T254 = T232[2'h3:2'h3];
  assign T255 = T241[1'h0:1'h0];
  assign T256 = T241[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T257 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T258 = state == 3'h1;
  assign io_outer_acquire_bits_union = T259;
  assign T259 = T258 ? oacq_probe_union : T260;
  assign T260 = T257 ? T267 : T261;
  assign T261 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T419;
  assign T419 = {4'h0, T262};
  assign T262 = {T263, 6'h0};
  assign T263 = {T266, T264};
  assign T264 = xact_union[4'h8:3'h6];
  assign T265 = T59 ? io_inner_acquire_bits_union : xact_union;
  assign T266 = xact_union[4'hc:4'h9];
  assign T267 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T268;
  assign T268 = {T269, 1'h1};
  assign T269 = 16'hffff;
  assign oacq_write_beat_union = T270;
  assign T270 = {T271, 1'h1};
  assign T271 = T288 ? T279 : T272;
  assign T272 = T274 ? T273 : 16'h0;
  assign T273 = xact_union[5'h10:1'h1];
  assign T274 = T277 | T275;
  assign T275 = xact_is_builtin_type & T276;
  assign T276 = xact_a_type == 3'h2;
  assign T277 = xact_is_builtin_type & T278;
  assign T278 = xact_a_type == 3'h3;
  assign T279 = T280;
  assign T280 = {T286, T281};
  assign T281 = 8'h0 - T420;
  assign T420 = {7'h0, T282};
  assign T282 = T283[1'h0:1'h0];
  assign T283 = 1'h1 << T284;
  assign T284 = T285[2'h3:2'h3];
  assign T285 = xact_union[4'hc:4'h9];
  assign T286 = 8'h0 - T421;
  assign T421 = {7'h0, T287};
  assign T287 = T283[1'h1:1'h1];
  assign T288 = xact_is_builtin_type & T289;
  assign T289 = xact_a_type == 3'h4;
  assign oacq_probe_union = T290;
  assign T290 = {T291, 1'h1};
  assign T291 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T292;
  assign T292 = T258 ? oacq_probe_a_type : T293;
  assign T293 = T257 ? T295 : T294;
  assign T294 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T295 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T296;
  assign T296 = T258 ? oacq_probe_is_builtin_type : T297;
  assign T297 = T257 ? T299 : T298;
  assign T298 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T299 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T300;
  assign T300 = T258 ? oacq_probe_addr_beat : T301;
  assign T301 = T257 ? T304 : T302;
  assign T302 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T303 = T59 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T304 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T305;
  assign T305 = T258 ? oacq_probe_client_xact_id : T306;
  assign T306 = T257 ? T308 : T307;
  assign T307 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h1;
  assign oacq_read_beat_client_xact_id = 4'h1;
  assign T308 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h1;
  assign oacq_write_beat_client_xact_id = 4'h1;
  assign oacq_probe_client_xact_id = 4'h1;
  assign io_outer_acquire_bits_addr_block = T309;
  assign T309 = T258 ? oacq_probe_addr_block : T310;
  assign T310 = T257 ? T312 : T311;
  assign T311 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T312 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T313;
  assign T313 = T124 ? T340 : T314;
  assign T314 = T121 ? T315 : T114;
  assign T315 = T339 & T316;
  assign T316 = T338 | T317;
  assign T317 = T322 & T318;
  assign T318 = T319 - 1'h1;
  assign T319 = 1'h1 << T320;
  assign T320 = T321 + 2'h1;
  assign T321 = oacq_data_cnt - oacq_data_cnt;
  assign T322 = iacq_data_valid >> oacq_data_cnt;
  assign T422 = reset ? 4'h0 : T323;
  assign T323 = T59 ? T331 : T324;
  assign T324 = T229 ? T325 : iacq_data_valid;
  assign T325 = T329 | T326;
  assign T326 = T423 & T327;
  assign T327 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T423 = T328 ? 4'hf : 4'h0;
  assign T328 = 1'h1;
  assign T329 = iacq_data_valid & T330;
  assign T330 = ~ T327;
  assign T331 = T332 << io_inner_acquire_bits_addr_beat;
  assign T332 = io_inner_acquire_bits_is_builtin_type & T333;
  assign T333 = T335 | T334;
  assign T334 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T335 = T337 | T336;
  assign T336 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T337 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T338 = collect_iacq_data ^ 1'h1;
  assign T339 = pending_ognt_ack ^ 1'h1;
  assign T340 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T341;
  assign T341 = T102 ? T342 : 1'h0;
  assign T342 = T343 | io_outer_acquire_ready;
  assign T343 = T344 ^ 1'h1;
  assign T344 = T346 | T345;
  assign T345 = 3'h2 == io_inner_release_bits_r_type;
  assign T346 = T348 | T347;
  assign T347 = 3'h1 == io_inner_release_bits_r_type;
  assign T348 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T349;
  assign T349 = T424;
  assign T424 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T356;
  assign T356 = T357;
  assign T357 = xact_is_builtin_type ? T362 : T358;
  assign T358 = T361 ? 2'h1 : T359;
  assign T359 = T360 ? 2'h0 : 2'h2;
  assign T360 = xact_a_type == 3'h1;
  assign T361 = xact_a_type == 3'h0;
  assign T362 = T371 ? 2'h2 : T363;
  assign T363 = T370 ? 2'h0 : T364;
  assign T364 = T369 ? 2'h2 : T365;
  assign T365 = T368 ? 2'h0 : T366;
  assign T366 = T367 ? 2'h0 : 2'h2;
  assign T367 = xact_a_type == 3'h4;
  assign T368 = xact_a_type == 3'h2;
  assign T369 = xact_a_type == 3'h0;
  assign T370 = xact_a_type == 3'h3;
  assign T371 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T372;
  assign T372 = xact_addr_block;
  assign io_inner_probe_valid = T373;
  assign T373 = T102 ? T374 : 1'h0;
  assign T374 = pending_probes != 1'h0;
  assign T425 = T426[1'h0:1'h0];
  assign T426 = reset ? 4'h0 : T350;
  assign T350 = T355 ? T428 : T351;
  assign T351 = T91 ? mask_incoherent : T427;
  assign T427 = {3'h0, pending_probes};
  assign T428 = {2'h0, T352};
  assign T352 = T429 & T353;
  assign T353 = ~ T354;
  assign T354 = 1'h1 << 1'h0;
  assign T429 = {1'h0, pending_probes};
  assign T355 = T102 & io_inner_probe_ready;
  assign io_inner_finish_ready = T150;
  assign io_inner_grant_bits_client_id = T375;
  assign T375 = xact_client_id;
  assign io_inner_grant_bits_data = T376;
  assign T376 = 4'h0;
  assign io_inner_grant_bits_g_type = T377;
  assign T377 = T430;
  assign T430 = {1'h0, T378};
  assign T378 = xact_is_builtin_type ? T381 : T431;
  assign T431 = {1'h0, T379};
  assign T379 = T380 ? 2'h0 : 2'h1;
  assign T380 = xact_a_type == 3'h0;
  assign T381 = T392 ? 3'h4 : T382;
  assign T382 = T391 ? 3'h5 : T383;
  assign T383 = T390 ? 3'h3 : T384;
  assign T384 = T389 ? 3'h3 : T385;
  assign T385 = T388 ? 3'h4 : T386;
  assign T386 = T387 ? 3'h1 : 3'h3;
  assign T387 = xact_a_type == 3'h5;
  assign T388 = xact_a_type == 3'h4;
  assign T389 = xact_a_type == 3'h3;
  assign T390 = xact_a_type == 3'h2;
  assign T391 = xact_a_type == 3'h1;
  assign T392 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T393;
  assign T393 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T394;
  assign T394 = 4'h1;
  assign io_inner_grant_bits_client_xact_id = T395;
  assign T395 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T396;
  assign T396 = 2'h0;
  assign io_inner_grant_valid = T397;
  assign T397 = T148 ? 1'h1 : T398;
  assign T398 = T142 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T399;
  assign T399 = T60 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T185 <= 1'b1;
  if(!T186 && T185 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T175 <= 1'b1;
  if(!T176 && T175 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T151 <= 1'b1;
  if(!T152 && T151 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= 3'h0;
    end else if(T147) begin
      state <= T143;
    end else if(T129) begin
      state <= T125;
    end else if(T122) begin
      state <= 3'h5;
    end else if(T120) begin
      state <= T119;
    end else if(T117) begin
      state <= T115;
    end else if(T76) begin
      state <= T61;
    end else if(T59) begin
      state <= T19;
    end
    if(T59) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T59) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T406;
    if(reset) begin
      R107 <= 2'h0;
    end else if(T110) begin
      R107 <= T109;
    end
    if(reset) begin
      R133 <= 2'h0;
    end else if(T136) begin
      R133 <= T135;
    end
    if(T59) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T59) begin
      collect_iacq_data <= T172;
    end else if(T162) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R166 <= 2'h0;
    end else if(T169) begin
      R166 <= T168;
    end
    if(T59) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T59) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T120) begin
      pending_ognt_ack <= 1'h1;
    end else if(T103) begin
      pending_ognt_ack <= 1'h1;
    end else if(T211) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T230) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T225) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T238) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T236) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T247) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T245) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T253) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T251) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T59) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T59) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T59) begin
      iacq_data_valid <= T331;
    end else if(T229) begin
      iacq_data_valid <= T325;
    end
    pending_probes <= T425;
  end
endmodule

module BroadcastAcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T400;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T401;
  wire[2:0] T25;
  wire[2:0] T402;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire pending_outer_write_;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[3:0] mask_incoherent;
  wire[3:0] T403;
  wire T51;
  wire T52;
  wire[3:0] mask_self;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T404;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T405;
  wire T58;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[2:0] T62;
  wire pending_outer_read;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire pending_outer_write;
  wire T69;
  wire T70;
  reg [2:0] xact_a_type;
  wire[2:0] T71;
  wire T72;
  wire T73;
  wire T74;
  reg  xact_is_builtin_type;
  wire T75;
  wire T76;
  wire T77;
  reg  release_count;
  wire T406;
  wire[2:0] T407;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T408;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire T85;
  wire[1:0] T409;
  wire T86;
  wire[2:0] T410;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T411;
  wire T90;
  wire T91;
  wire[2:0] T412;
  wire T92;
  wire[2:0] T413;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire oacq_data_done;
  wire T104;
  wire T105;
  wire T106;
  reg [1:0] R107;
  wire[1:0] T414;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire[2:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire ignt_data_done;
  wire T130;
  wire T131;
  wire T132;
  reg [1:0] R133;
  wire[1:0] T415;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire[2:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  reg[0:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire T159;
  reg  collect_iacq_data;
  wire T416;
  wire T160;
  wire T161;
  wire T162;
  wire iacq_data_done;
  wire T163;
  wire T164;
  wire T165;
  reg [1:0] R166;
  wire[1:0] T417;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  reg[0:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  reg [1:0] xact_client_id;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  reg[0:0] T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  reg [25:0] xact_addr_block;
  wire[25:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  reg  pending_ognt_ack;
  wire T418;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[3:0] T214;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[3:0] T220;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T221;
  wire[3:0] T222;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T223;
  wire[3:0] T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[1:0] T228;
  wire T229;
  wire T230;
  wire T231;
  wire[3:0] T232;
  wire[1:0] T233;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T234;
  wire[3:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[1:0] T241;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T242;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T243;
  wire[3:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T249;
  wire[3:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] oacq_write_beat_data;
  wire T257;
  wire[3:0] oacq_probe_data;
  wire T258;
  wire[16:0] T259;
  wire[16:0] T260;
  wire[16:0] T261;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T419;
  wire[12:0] T262;
  wire[6:0] T263;
  wire[2:0] T264;
  reg [16:0] xact_union;
  wire[16:0] T265;
  wire[3:0] T266;
  wire[16:0] T267;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T268;
  wire[15:0] T269;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T270;
  wire[15:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[15:0] T279;
  wire[15:0] T280;
  wire[7:0] T281;
  wire[7:0] T420;
  wire T282;
  wire[1:0] T283;
  wire T284;
  wire[3:0] T285;
  wire[7:0] T286;
  wire[7:0] T421;
  wire T287;
  wire T288;
  wire T289;
  wire[16:0] oacq_probe_union;
  wire[16:0] T290;
  wire[15:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[2:0] T294;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T295;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T296;
  wire T297;
  wire T298;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T299;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T303;
  wire[1:0] T304;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T308;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T309;
  wire[25:0] T310;
  wire[25:0] T311;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T312;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire[1:0] T321;
  wire T322;
  reg [3:0] iacq_data_valid;
  wire[3:0] T422;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[3:0] T326;
  wire[3:0] T327;
  wire[3:0] T423;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire[1:0] T349;
  wire[1:0] T424;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[1:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[25:0] T372;
  wire T373;
  wire T374;
  reg  pending_probes;
  wire T425;
  wire[3:0] T426;
  wire[3:0] T350;
  wire[3:0] T351;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[1:0] T352;
  wire T353;
  wire T354;
  wire[1:0] T429;
  wire T355;
  wire[1:0] T375;
  wire[3:0] T376;
  wire[3:0] T377;
  wire[3:0] T430;
  wire[2:0] T378;
  wire[2:0] T431;
  wire[1:0] T379;
  wire T380;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] T384;
  wire[2:0] T385;
  wire[2:0] T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[3:0] T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire T397;
  wire T398;
  wire T399;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R107 = {1{$random}};
    R133 = {1{$random}};
    T151 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R166 = {1{$random}};
    T175 = 1'b0;
    xact_client_id = {1{$random}};
    T185 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T400 = reset ? 3'h0 : T11;
  assign T11 = T149 ? 3'h0 : T12;
  assign T12 = T147 ? T143 : T13;
  assign T13 = T129 ? T125 : T14;
  assign T14 = T122 ? 3'h5 : T15;
  assign T15 = T120 ? T119 : T16;
  assign T16 = T117 ? T115 : T17;
  assign T17 = T76 ? T61 : T18;
  assign T18 = T59 ? T19 : state;
  assign T19 = T50 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T44 ? T41 : T22;
  assign T22 = T40 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T401;
  assign T401 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T402;
  assign T402 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T39 ? 3'h4 : T29;
  assign T29 = T38 ? 3'h5 : T30;
  assign T30 = T37 ? 3'h3 : T31;
  assign T31 = T36 ? 3'h3 : T32;
  assign T32 = T35 ? 3'h4 : T33;
  assign T33 = T34 ? 3'h1 : 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h5;
  assign T35 = io_inner_acquire_bits_a_type == 3'h4;
  assign T36 = io_inner_acquire_bits_a_type == 3'h3;
  assign T37 = io_inner_acquire_bits_a_type == 3'h2;
  assign T38 = io_inner_acquire_bits_a_type == 3'h1;
  assign T39 = io_inner_acquire_bits_a_type == 3'h0;
  assign T40 = 4'h0 == T24;
  assign T41 = T43 | T42;
  assign T42 = 4'h4 == T24;
  assign T43 = 4'h5 == T24;
  assign T44 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T45;
  assign T45 = T47 | T46;
  assign T46 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T49 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T50 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T403;
  assign T403 = {3'h0, T51};
  assign T51 = ~ T52;
  assign T52 = io_incoherent_0;
  assign mask_self = T56 | T53;
  assign T53 = T404 & T54;
  assign T54 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T404 = T55 ? 4'hf : 4'h0;
  assign T55 = 1'h0;
  assign T56 = T405 & T57;
  assign T57 = ~ T54;
  assign T405 = {3'h0, T58};
  assign T58 = 1'h1;
  assign T59 = T60 & io_inner_acquire_valid;
  assign T60 = 3'h0 == state;
  assign T61 = pending_outer_write ? 3'h3 : T62;
  assign T62 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T66 : T63;
  assign T63 = T65 | T64;
  assign T64 = 4'h1 == io_inner_grant_bits_g_type;
  assign T65 = 4'h0 == io_inner_grant_bits_g_type;
  assign T66 = T68 | T67;
  assign T67 = 4'h4 == io_inner_grant_bits_g_type;
  assign T68 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T69;
  assign T69 = T72 | T70;
  assign T70 = 3'h4 == xact_a_type;
  assign T71 = T59 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T72 = T74 | T73;
  assign T73 = 3'h3 == xact_a_type;
  assign T74 = 3'h2 == xact_a_type;
  assign T75 = T59 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T76 = T103 & T77;
  assign T77 = release_count == 1'h1;
  assign T406 = T407[1'h0:1'h0];
  assign T407 = reset ? 3'h0 : T78;
  assign T78 = T94 ? T413 : T79;
  assign T79 = T103 ? T412 : T80;
  assign T80 = T91 ? T81 : T408;
  assign T408 = {2'h0, release_count};
  assign T81 = T410 + T82;
  assign T82 = {1'h0, T83};
  assign T83 = T409 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = mask_incoherent[2'h3:2'h3];
  assign T409 = {1'h0, T86};
  assign T86 = mask_incoherent[2'h2:2'h2];
  assign T410 = {1'h0, T87};
  assign T87 = T411 + T88;
  assign T88 = {1'h0, T89};
  assign T89 = mask_incoherent[1'h1:1'h1];
  assign T411 = {1'h0, T90};
  assign T90 = mask_incoherent[1'h0:1'h0];
  assign T91 = T59 & T50;
  assign T412 = {2'h0, T92};
  assign T92 = release_count - 1'h1;
  assign T413 = {2'h0, T93};
  assign T93 = release_count - 1'h1;
  assign T94 = T101 & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = T98 | T97;
  assign T97 = 3'h2 == io_inner_release_bits_r_type;
  assign T98 = T100 | T99;
  assign T99 = 3'h1 == io_inner_release_bits_r_type;
  assign T100 = 3'h0 == io_inner_release_bits_r_type;
  assign T101 = T102 & io_inner_release_valid;
  assign T102 = 3'h1 == state;
  assign T103 = T113 & oacq_data_done;
  assign oacq_data_done = T111 ? T105 : T104;
  assign T104 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T105 = T110 & T106;
  assign T106 = R107 == 2'h3;
  assign T414 = reset ? 2'h0 : T108;
  assign T108 = T110 ? T109 : R107;
  assign T109 = R107 + 2'h1;
  assign T110 = T104 & T111;
  assign T111 = io_outer_acquire_bits_is_builtin_type & T112;
  assign T112 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T113 = T114 & io_outer_acquire_ready;
  assign T114 = T101 & T96;
  assign T115 = pending_outer_write ? 3'h3 : T116;
  assign T116 = pending_outer_read ? 3'h2 : 3'h4;
  assign T117 = T94 & T118;
  assign T118 = release_count == 1'h1;
  assign T119 = pending_outer_read ? 3'h2 : 3'h5;
  assign T120 = T121 & oacq_data_done;
  assign T121 = 3'h3 == state;
  assign T122 = T124 & T123;
  assign T123 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T124 = 3'h2 == state;
  assign T125 = T126 ? 3'h6 : 3'h0;
  assign T126 = T127 ^ 1'h1;
  assign T127 = io_inner_grant_bits_is_builtin_type & T128;
  assign T128 = io_inner_grant_bits_g_type == 4'h0;
  assign T129 = T142 & ignt_data_done;
  assign ignt_data_done = T137 ? T131 : T130;
  assign T130 = io_inner_grant_ready & io_inner_grant_valid;
  assign T131 = T136 & T132;
  assign T132 = R133 == 2'h3;
  assign T415 = reset ? 2'h0 : T134;
  assign T134 = T136 ? T135 : R133;
  assign T135 = R133 + 2'h1;
  assign T136 = T130 & T137;
  assign T137 = io_inner_grant_bits_is_builtin_type ? T141 : T138;
  assign T138 = T140 | T139;
  assign T139 = 4'h1 == io_inner_grant_bits_g_type;
  assign T140 = 4'h0 == io_inner_grant_bits_g_type;
  assign T141 = 4'h5 == io_inner_grant_bits_g_type;
  assign T142 = 3'h5 == state;
  assign T143 = T144 ? 3'h6 : 3'h0;
  assign T144 = T145 ^ 1'h1;
  assign T145 = io_inner_grant_bits_is_builtin_type & T146;
  assign T146 = io_inner_grant_bits_g_type == 4'h0;
  assign T147 = T148 & io_inner_grant_ready;
  assign T148 = 3'h4 == state;
  assign T149 = T150 & io_inner_finish_valid;
  assign T150 = 3'h6 == state;
  assign T152 = T153 | reset;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T157 & T155;
  assign T155 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T156 = T59 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T157 = T159 & T158;
  assign T158 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T159 = T174 & collect_iacq_data;
  assign T416 = reset ? 1'h0 : T160;
  assign T160 = T59 ? T172 : T161;
  assign T161 = T162 ? 1'h0 : collect_iacq_data;
  assign T162 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T170 ? T164 : T163;
  assign T163 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T164 = T169 & T165;
  assign T165 = R166 == 2'h3;
  assign T417 = reset ? 2'h0 : T167;
  assign T167 = T169 ? T168 : R166;
  assign T168 = R166 + 2'h1;
  assign T169 = T163 & T170;
  assign T170 = io_inner_acquire_bits_is_builtin_type & T171;
  assign T171 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = state != 3'h0;
  assign T176 = T177 | reset;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T181 & T179;
  assign T179 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T180 = T59 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T181 = T183 & T182;
  assign T182 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T183 = T184 & collect_iacq_data;
  assign T184 = state != 3'h0;
  assign T186 = T187 | reset;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T192 & T189;
  assign T189 = T191 | T190;
  assign T190 = 3'h5 == xact_a_type;
  assign T191 = 3'h4 == xact_a_type;
  assign T192 = T193 & xact_is_builtin_type;
  assign T193 = state != 3'h0;
  assign io_has_release_match = T194;
  assign T194 = T196 & T195;
  assign T195 = state == 3'h1;
  assign T196 = T198 & T197;
  assign T197 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T198 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T199 = T59 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T200;
  assign T200 = T201 & collect_iacq_data;
  assign T201 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T202;
  assign T202 = T204 & T203;
  assign T203 = collect_iacq_data ^ 1'h1;
  assign T204 = T206 & T205;
  assign T205 = state != 3'h0;
  assign T206 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T207;
  assign T207 = T142 ? io_inner_grant_ready : pending_ognt_ack;
  assign T418 = reset ? 1'h0 : T208;
  assign T208 = T120 ? 1'h1 : T209;
  assign T209 = T103 ? 1'h1 : T210;
  assign T210 = T211 ? 1'h0 : pending_ognt_ack;
  assign T211 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T212;
  assign T212 = T258 ? oacq_probe_data : T213;
  assign T213 = T257 ? T220 : T214;
  assign T214 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T215;
  assign T215 = T217 | T216;
  assign T216 = 3'h4 == xact_a_type;
  assign T217 = T219 | T218;
  assign T218 = 3'h0 == xact_a_type;
  assign T219 = 3'h2 == xact_a_type;
  assign T220 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T221;
  assign T221 = T256 ? T242 : T222;
  assign T222 = T240 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T223 = T230 ? io_inner_acquire_bits_data : T224;
  assign T224 = T225 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T225 = T229 & T226;
  assign T226 = T227[1'h0:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = io_inner_acquire_bits_addr_beat;
  assign T229 = collect_iacq_data & io_inner_acquire_valid;
  assign T230 = T59 & T231;
  assign T231 = T232[1'h0:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = 2'h0;
  assign T234 = T238 ? io_inner_acquire_bits_data : T235;
  assign T235 = T236 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T236 = T229 & T237;
  assign T237 = T227[1'h1:1'h1];
  assign T238 = T59 & T239;
  assign T239 = T232[1'h1:1'h1];
  assign T240 = T241[1'h0:1'h0];
  assign T241 = oacq_data_cnt;
  assign oacq_data_cnt = T111 ? R107 : 2'h0;
  assign T242 = T255 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T243 = T247 ? io_inner_acquire_bits_data : T244;
  assign T244 = T245 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T245 = T229 & T246;
  assign T246 = T227[2'h2:2'h2];
  assign T247 = T59 & T248;
  assign T248 = T232[2'h2:2'h2];
  assign T249 = T253 ? io_inner_acquire_bits_data : T250;
  assign T250 = T251 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T251 = T229 & T252;
  assign T252 = T227[2'h3:2'h3];
  assign T253 = T59 & T254;
  assign T254 = T232[2'h3:2'h3];
  assign T255 = T241[1'h0:1'h0];
  assign T256 = T241[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T257 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T258 = state == 3'h1;
  assign io_outer_acquire_bits_union = T259;
  assign T259 = T258 ? oacq_probe_union : T260;
  assign T260 = T257 ? T267 : T261;
  assign T261 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T419;
  assign T419 = {4'h0, T262};
  assign T262 = {T263, 6'h0};
  assign T263 = {T266, T264};
  assign T264 = xact_union[4'h8:3'h6];
  assign T265 = T59 ? io_inner_acquire_bits_union : xact_union;
  assign T266 = xact_union[4'hc:4'h9];
  assign T267 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T268;
  assign T268 = {T269, 1'h1};
  assign T269 = 16'hffff;
  assign oacq_write_beat_union = T270;
  assign T270 = {T271, 1'h1};
  assign T271 = T288 ? T279 : T272;
  assign T272 = T274 ? T273 : 16'h0;
  assign T273 = xact_union[5'h10:1'h1];
  assign T274 = T277 | T275;
  assign T275 = xact_is_builtin_type & T276;
  assign T276 = xact_a_type == 3'h2;
  assign T277 = xact_is_builtin_type & T278;
  assign T278 = xact_a_type == 3'h3;
  assign T279 = T280;
  assign T280 = {T286, T281};
  assign T281 = 8'h0 - T420;
  assign T420 = {7'h0, T282};
  assign T282 = T283[1'h0:1'h0];
  assign T283 = 1'h1 << T284;
  assign T284 = T285[2'h3:2'h3];
  assign T285 = xact_union[4'hc:4'h9];
  assign T286 = 8'h0 - T421;
  assign T421 = {7'h0, T287};
  assign T287 = T283[1'h1:1'h1];
  assign T288 = xact_is_builtin_type & T289;
  assign T289 = xact_a_type == 3'h4;
  assign oacq_probe_union = T290;
  assign T290 = {T291, 1'h1};
  assign T291 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T292;
  assign T292 = T258 ? oacq_probe_a_type : T293;
  assign T293 = T257 ? T295 : T294;
  assign T294 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T295 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T296;
  assign T296 = T258 ? oacq_probe_is_builtin_type : T297;
  assign T297 = T257 ? T299 : T298;
  assign T298 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T299 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T300;
  assign T300 = T258 ? oacq_probe_addr_beat : T301;
  assign T301 = T257 ? T304 : T302;
  assign T302 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T303 = T59 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T304 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T305;
  assign T305 = T258 ? oacq_probe_client_xact_id : T306;
  assign T306 = T257 ? T308 : T307;
  assign T307 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h2;
  assign oacq_read_beat_client_xact_id = 4'h2;
  assign T308 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h2;
  assign oacq_write_beat_client_xact_id = 4'h2;
  assign oacq_probe_client_xact_id = 4'h2;
  assign io_outer_acquire_bits_addr_block = T309;
  assign T309 = T258 ? oacq_probe_addr_block : T310;
  assign T310 = T257 ? T312 : T311;
  assign T311 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T312 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T313;
  assign T313 = T124 ? T340 : T314;
  assign T314 = T121 ? T315 : T114;
  assign T315 = T339 & T316;
  assign T316 = T338 | T317;
  assign T317 = T322 & T318;
  assign T318 = T319 - 1'h1;
  assign T319 = 1'h1 << T320;
  assign T320 = T321 + 2'h1;
  assign T321 = oacq_data_cnt - oacq_data_cnt;
  assign T322 = iacq_data_valid >> oacq_data_cnt;
  assign T422 = reset ? 4'h0 : T323;
  assign T323 = T59 ? T331 : T324;
  assign T324 = T229 ? T325 : iacq_data_valid;
  assign T325 = T329 | T326;
  assign T326 = T423 & T327;
  assign T327 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T423 = T328 ? 4'hf : 4'h0;
  assign T328 = 1'h1;
  assign T329 = iacq_data_valid & T330;
  assign T330 = ~ T327;
  assign T331 = T332 << io_inner_acquire_bits_addr_beat;
  assign T332 = io_inner_acquire_bits_is_builtin_type & T333;
  assign T333 = T335 | T334;
  assign T334 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T335 = T337 | T336;
  assign T336 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T337 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T338 = collect_iacq_data ^ 1'h1;
  assign T339 = pending_ognt_ack ^ 1'h1;
  assign T340 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T341;
  assign T341 = T102 ? T342 : 1'h0;
  assign T342 = T343 | io_outer_acquire_ready;
  assign T343 = T344 ^ 1'h1;
  assign T344 = T346 | T345;
  assign T345 = 3'h2 == io_inner_release_bits_r_type;
  assign T346 = T348 | T347;
  assign T347 = 3'h1 == io_inner_release_bits_r_type;
  assign T348 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T349;
  assign T349 = T424;
  assign T424 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T356;
  assign T356 = T357;
  assign T357 = xact_is_builtin_type ? T362 : T358;
  assign T358 = T361 ? 2'h1 : T359;
  assign T359 = T360 ? 2'h0 : 2'h2;
  assign T360 = xact_a_type == 3'h1;
  assign T361 = xact_a_type == 3'h0;
  assign T362 = T371 ? 2'h2 : T363;
  assign T363 = T370 ? 2'h0 : T364;
  assign T364 = T369 ? 2'h2 : T365;
  assign T365 = T368 ? 2'h0 : T366;
  assign T366 = T367 ? 2'h0 : 2'h2;
  assign T367 = xact_a_type == 3'h4;
  assign T368 = xact_a_type == 3'h2;
  assign T369 = xact_a_type == 3'h0;
  assign T370 = xact_a_type == 3'h3;
  assign T371 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T372;
  assign T372 = xact_addr_block;
  assign io_inner_probe_valid = T373;
  assign T373 = T102 ? T374 : 1'h0;
  assign T374 = pending_probes != 1'h0;
  assign T425 = T426[1'h0:1'h0];
  assign T426 = reset ? 4'h0 : T350;
  assign T350 = T355 ? T428 : T351;
  assign T351 = T91 ? mask_incoherent : T427;
  assign T427 = {3'h0, pending_probes};
  assign T428 = {2'h0, T352};
  assign T352 = T429 & T353;
  assign T353 = ~ T354;
  assign T354 = 1'h1 << 1'h0;
  assign T429 = {1'h0, pending_probes};
  assign T355 = T102 & io_inner_probe_ready;
  assign io_inner_finish_ready = T150;
  assign io_inner_grant_bits_client_id = T375;
  assign T375 = xact_client_id;
  assign io_inner_grant_bits_data = T376;
  assign T376 = 4'h0;
  assign io_inner_grant_bits_g_type = T377;
  assign T377 = T430;
  assign T430 = {1'h0, T378};
  assign T378 = xact_is_builtin_type ? T381 : T431;
  assign T431 = {1'h0, T379};
  assign T379 = T380 ? 2'h0 : 2'h1;
  assign T380 = xact_a_type == 3'h0;
  assign T381 = T392 ? 3'h4 : T382;
  assign T382 = T391 ? 3'h5 : T383;
  assign T383 = T390 ? 3'h3 : T384;
  assign T384 = T389 ? 3'h3 : T385;
  assign T385 = T388 ? 3'h4 : T386;
  assign T386 = T387 ? 3'h1 : 3'h3;
  assign T387 = xact_a_type == 3'h5;
  assign T388 = xact_a_type == 3'h4;
  assign T389 = xact_a_type == 3'h3;
  assign T390 = xact_a_type == 3'h2;
  assign T391 = xact_a_type == 3'h1;
  assign T392 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T393;
  assign T393 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T394;
  assign T394 = 4'h2;
  assign io_inner_grant_bits_client_xact_id = T395;
  assign T395 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T396;
  assign T396 = 2'h0;
  assign io_inner_grant_valid = T397;
  assign T397 = T148 ? 1'h1 : T398;
  assign T398 = T142 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T399;
  assign T399 = T60 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T185 <= 1'b1;
  if(!T186 && T185 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T175 <= 1'b1;
  if(!T176 && T175 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T151 <= 1'b1;
  if(!T152 && T151 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= 3'h0;
    end else if(T147) begin
      state <= T143;
    end else if(T129) begin
      state <= T125;
    end else if(T122) begin
      state <= 3'h5;
    end else if(T120) begin
      state <= T119;
    end else if(T117) begin
      state <= T115;
    end else if(T76) begin
      state <= T61;
    end else if(T59) begin
      state <= T19;
    end
    if(T59) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T59) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T406;
    if(reset) begin
      R107 <= 2'h0;
    end else if(T110) begin
      R107 <= T109;
    end
    if(reset) begin
      R133 <= 2'h0;
    end else if(T136) begin
      R133 <= T135;
    end
    if(T59) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T59) begin
      collect_iacq_data <= T172;
    end else if(T162) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R166 <= 2'h0;
    end else if(T169) begin
      R166 <= T168;
    end
    if(T59) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T59) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T120) begin
      pending_ognt_ack <= 1'h1;
    end else if(T103) begin
      pending_ognt_ack <= 1'h1;
    end else if(T211) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T230) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T225) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T238) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T236) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T247) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T245) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T253) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T251) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T59) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T59) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T59) begin
      iacq_data_valid <= T331;
    end else if(T229) begin
      iacq_data_valid <= T325;
    end
    pending_probes <= T425;
  end
endmodule

module BroadcastAcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T400;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T401;
  wire[2:0] T25;
  wire[2:0] T402;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire pending_outer_write_;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[3:0] mask_incoherent;
  wire[3:0] T403;
  wire T51;
  wire T52;
  wire[3:0] mask_self;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T404;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T405;
  wire T58;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[2:0] T62;
  wire pending_outer_read;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire pending_outer_write;
  wire T69;
  wire T70;
  reg [2:0] xact_a_type;
  wire[2:0] T71;
  wire T72;
  wire T73;
  wire T74;
  reg  xact_is_builtin_type;
  wire T75;
  wire T76;
  wire T77;
  reg  release_count;
  wire T406;
  wire[2:0] T407;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T408;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire T85;
  wire[1:0] T409;
  wire T86;
  wire[2:0] T410;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T411;
  wire T90;
  wire T91;
  wire[2:0] T412;
  wire T92;
  wire[2:0] T413;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire oacq_data_done;
  wire T104;
  wire T105;
  wire T106;
  reg [1:0] R107;
  wire[1:0] T414;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire[2:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire ignt_data_done;
  wire T130;
  wire T131;
  wire T132;
  reg [1:0] R133;
  wire[1:0] T415;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire[2:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  reg[0:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire T159;
  reg  collect_iacq_data;
  wire T416;
  wire T160;
  wire T161;
  wire T162;
  wire iacq_data_done;
  wire T163;
  wire T164;
  wire T165;
  reg [1:0] R166;
  wire[1:0] T417;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  reg[0:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  reg [1:0] xact_client_id;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  reg[0:0] T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  reg [25:0] xact_addr_block;
  wire[25:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  reg  pending_ognt_ack;
  wire T418;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[3:0] T214;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[3:0] T220;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T221;
  wire[3:0] T222;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T223;
  wire[3:0] T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[1:0] T228;
  wire T229;
  wire T230;
  wire T231;
  wire[3:0] T232;
  wire[1:0] T233;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T234;
  wire[3:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[1:0] T241;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T242;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T243;
  wire[3:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T249;
  wire[3:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] oacq_write_beat_data;
  wire T257;
  wire[3:0] oacq_probe_data;
  wire T258;
  wire[16:0] T259;
  wire[16:0] T260;
  wire[16:0] T261;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T419;
  wire[12:0] T262;
  wire[6:0] T263;
  wire[2:0] T264;
  reg [16:0] xact_union;
  wire[16:0] T265;
  wire[3:0] T266;
  wire[16:0] T267;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T268;
  wire[15:0] T269;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T270;
  wire[15:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[15:0] T279;
  wire[15:0] T280;
  wire[7:0] T281;
  wire[7:0] T420;
  wire T282;
  wire[1:0] T283;
  wire T284;
  wire[3:0] T285;
  wire[7:0] T286;
  wire[7:0] T421;
  wire T287;
  wire T288;
  wire T289;
  wire[16:0] oacq_probe_union;
  wire[16:0] T290;
  wire[15:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[2:0] T294;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T295;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T296;
  wire T297;
  wire T298;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T299;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T303;
  wire[1:0] T304;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T308;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T309;
  wire[25:0] T310;
  wire[25:0] T311;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T312;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire[1:0] T321;
  wire T322;
  reg [3:0] iacq_data_valid;
  wire[3:0] T422;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[3:0] T326;
  wire[3:0] T327;
  wire[3:0] T423;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire[1:0] T349;
  wire[1:0] T424;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[1:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[25:0] T372;
  wire T373;
  wire T374;
  reg  pending_probes;
  wire T425;
  wire[3:0] T426;
  wire[3:0] T350;
  wire[3:0] T351;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[1:0] T352;
  wire T353;
  wire T354;
  wire[1:0] T429;
  wire T355;
  wire[1:0] T375;
  wire[3:0] T376;
  wire[3:0] T377;
  wire[3:0] T430;
  wire[2:0] T378;
  wire[2:0] T431;
  wire[1:0] T379;
  wire T380;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] T384;
  wire[2:0] T385;
  wire[2:0] T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[3:0] T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire T397;
  wire T398;
  wire T399;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R107 = {1{$random}};
    R133 = {1{$random}};
    T151 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R166 = {1{$random}};
    T175 = 1'b0;
    xact_client_id = {1{$random}};
    T185 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T400 = reset ? 3'h0 : T11;
  assign T11 = T149 ? 3'h0 : T12;
  assign T12 = T147 ? T143 : T13;
  assign T13 = T129 ? T125 : T14;
  assign T14 = T122 ? 3'h5 : T15;
  assign T15 = T120 ? T119 : T16;
  assign T16 = T117 ? T115 : T17;
  assign T17 = T76 ? T61 : T18;
  assign T18 = T59 ? T19 : state;
  assign T19 = T50 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T44 ? T41 : T22;
  assign T22 = T40 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T401;
  assign T401 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T402;
  assign T402 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T39 ? 3'h4 : T29;
  assign T29 = T38 ? 3'h5 : T30;
  assign T30 = T37 ? 3'h3 : T31;
  assign T31 = T36 ? 3'h3 : T32;
  assign T32 = T35 ? 3'h4 : T33;
  assign T33 = T34 ? 3'h1 : 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h5;
  assign T35 = io_inner_acquire_bits_a_type == 3'h4;
  assign T36 = io_inner_acquire_bits_a_type == 3'h3;
  assign T37 = io_inner_acquire_bits_a_type == 3'h2;
  assign T38 = io_inner_acquire_bits_a_type == 3'h1;
  assign T39 = io_inner_acquire_bits_a_type == 3'h0;
  assign T40 = 4'h0 == T24;
  assign T41 = T43 | T42;
  assign T42 = 4'h4 == T24;
  assign T43 = 4'h5 == T24;
  assign T44 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T45;
  assign T45 = T47 | T46;
  assign T46 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T49 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T50 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T403;
  assign T403 = {3'h0, T51};
  assign T51 = ~ T52;
  assign T52 = io_incoherent_0;
  assign mask_self = T56 | T53;
  assign T53 = T404 & T54;
  assign T54 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T404 = T55 ? 4'hf : 4'h0;
  assign T55 = 1'h0;
  assign T56 = T405 & T57;
  assign T57 = ~ T54;
  assign T405 = {3'h0, T58};
  assign T58 = 1'h1;
  assign T59 = T60 & io_inner_acquire_valid;
  assign T60 = 3'h0 == state;
  assign T61 = pending_outer_write ? 3'h3 : T62;
  assign T62 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T66 : T63;
  assign T63 = T65 | T64;
  assign T64 = 4'h1 == io_inner_grant_bits_g_type;
  assign T65 = 4'h0 == io_inner_grant_bits_g_type;
  assign T66 = T68 | T67;
  assign T67 = 4'h4 == io_inner_grant_bits_g_type;
  assign T68 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T69;
  assign T69 = T72 | T70;
  assign T70 = 3'h4 == xact_a_type;
  assign T71 = T59 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T72 = T74 | T73;
  assign T73 = 3'h3 == xact_a_type;
  assign T74 = 3'h2 == xact_a_type;
  assign T75 = T59 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T76 = T103 & T77;
  assign T77 = release_count == 1'h1;
  assign T406 = T407[1'h0:1'h0];
  assign T407 = reset ? 3'h0 : T78;
  assign T78 = T94 ? T413 : T79;
  assign T79 = T103 ? T412 : T80;
  assign T80 = T91 ? T81 : T408;
  assign T408 = {2'h0, release_count};
  assign T81 = T410 + T82;
  assign T82 = {1'h0, T83};
  assign T83 = T409 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = mask_incoherent[2'h3:2'h3];
  assign T409 = {1'h0, T86};
  assign T86 = mask_incoherent[2'h2:2'h2];
  assign T410 = {1'h0, T87};
  assign T87 = T411 + T88;
  assign T88 = {1'h0, T89};
  assign T89 = mask_incoherent[1'h1:1'h1];
  assign T411 = {1'h0, T90};
  assign T90 = mask_incoherent[1'h0:1'h0];
  assign T91 = T59 & T50;
  assign T412 = {2'h0, T92};
  assign T92 = release_count - 1'h1;
  assign T413 = {2'h0, T93};
  assign T93 = release_count - 1'h1;
  assign T94 = T101 & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = T98 | T97;
  assign T97 = 3'h2 == io_inner_release_bits_r_type;
  assign T98 = T100 | T99;
  assign T99 = 3'h1 == io_inner_release_bits_r_type;
  assign T100 = 3'h0 == io_inner_release_bits_r_type;
  assign T101 = T102 & io_inner_release_valid;
  assign T102 = 3'h1 == state;
  assign T103 = T113 & oacq_data_done;
  assign oacq_data_done = T111 ? T105 : T104;
  assign T104 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T105 = T110 & T106;
  assign T106 = R107 == 2'h3;
  assign T414 = reset ? 2'h0 : T108;
  assign T108 = T110 ? T109 : R107;
  assign T109 = R107 + 2'h1;
  assign T110 = T104 & T111;
  assign T111 = io_outer_acquire_bits_is_builtin_type & T112;
  assign T112 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T113 = T114 & io_outer_acquire_ready;
  assign T114 = T101 & T96;
  assign T115 = pending_outer_write ? 3'h3 : T116;
  assign T116 = pending_outer_read ? 3'h2 : 3'h4;
  assign T117 = T94 & T118;
  assign T118 = release_count == 1'h1;
  assign T119 = pending_outer_read ? 3'h2 : 3'h5;
  assign T120 = T121 & oacq_data_done;
  assign T121 = 3'h3 == state;
  assign T122 = T124 & T123;
  assign T123 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T124 = 3'h2 == state;
  assign T125 = T126 ? 3'h6 : 3'h0;
  assign T126 = T127 ^ 1'h1;
  assign T127 = io_inner_grant_bits_is_builtin_type & T128;
  assign T128 = io_inner_grant_bits_g_type == 4'h0;
  assign T129 = T142 & ignt_data_done;
  assign ignt_data_done = T137 ? T131 : T130;
  assign T130 = io_inner_grant_ready & io_inner_grant_valid;
  assign T131 = T136 & T132;
  assign T132 = R133 == 2'h3;
  assign T415 = reset ? 2'h0 : T134;
  assign T134 = T136 ? T135 : R133;
  assign T135 = R133 + 2'h1;
  assign T136 = T130 & T137;
  assign T137 = io_inner_grant_bits_is_builtin_type ? T141 : T138;
  assign T138 = T140 | T139;
  assign T139 = 4'h1 == io_inner_grant_bits_g_type;
  assign T140 = 4'h0 == io_inner_grant_bits_g_type;
  assign T141 = 4'h5 == io_inner_grant_bits_g_type;
  assign T142 = 3'h5 == state;
  assign T143 = T144 ? 3'h6 : 3'h0;
  assign T144 = T145 ^ 1'h1;
  assign T145 = io_inner_grant_bits_is_builtin_type & T146;
  assign T146 = io_inner_grant_bits_g_type == 4'h0;
  assign T147 = T148 & io_inner_grant_ready;
  assign T148 = 3'h4 == state;
  assign T149 = T150 & io_inner_finish_valid;
  assign T150 = 3'h6 == state;
  assign T152 = T153 | reset;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T157 & T155;
  assign T155 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T156 = T59 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T157 = T159 & T158;
  assign T158 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T159 = T174 & collect_iacq_data;
  assign T416 = reset ? 1'h0 : T160;
  assign T160 = T59 ? T172 : T161;
  assign T161 = T162 ? 1'h0 : collect_iacq_data;
  assign T162 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T170 ? T164 : T163;
  assign T163 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T164 = T169 & T165;
  assign T165 = R166 == 2'h3;
  assign T417 = reset ? 2'h0 : T167;
  assign T167 = T169 ? T168 : R166;
  assign T168 = R166 + 2'h1;
  assign T169 = T163 & T170;
  assign T170 = io_inner_acquire_bits_is_builtin_type & T171;
  assign T171 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = state != 3'h0;
  assign T176 = T177 | reset;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T181 & T179;
  assign T179 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T180 = T59 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T181 = T183 & T182;
  assign T182 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T183 = T184 & collect_iacq_data;
  assign T184 = state != 3'h0;
  assign T186 = T187 | reset;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T192 & T189;
  assign T189 = T191 | T190;
  assign T190 = 3'h5 == xact_a_type;
  assign T191 = 3'h4 == xact_a_type;
  assign T192 = T193 & xact_is_builtin_type;
  assign T193 = state != 3'h0;
  assign io_has_release_match = T194;
  assign T194 = T196 & T195;
  assign T195 = state == 3'h1;
  assign T196 = T198 & T197;
  assign T197 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T198 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T199 = T59 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T200;
  assign T200 = T201 & collect_iacq_data;
  assign T201 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T202;
  assign T202 = T204 & T203;
  assign T203 = collect_iacq_data ^ 1'h1;
  assign T204 = T206 & T205;
  assign T205 = state != 3'h0;
  assign T206 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T207;
  assign T207 = T142 ? io_inner_grant_ready : pending_ognt_ack;
  assign T418 = reset ? 1'h0 : T208;
  assign T208 = T120 ? 1'h1 : T209;
  assign T209 = T103 ? 1'h1 : T210;
  assign T210 = T211 ? 1'h0 : pending_ognt_ack;
  assign T211 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T212;
  assign T212 = T258 ? oacq_probe_data : T213;
  assign T213 = T257 ? T220 : T214;
  assign T214 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T215;
  assign T215 = T217 | T216;
  assign T216 = 3'h4 == xact_a_type;
  assign T217 = T219 | T218;
  assign T218 = 3'h0 == xact_a_type;
  assign T219 = 3'h2 == xact_a_type;
  assign T220 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T221;
  assign T221 = T256 ? T242 : T222;
  assign T222 = T240 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T223 = T230 ? io_inner_acquire_bits_data : T224;
  assign T224 = T225 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T225 = T229 & T226;
  assign T226 = T227[1'h0:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = io_inner_acquire_bits_addr_beat;
  assign T229 = collect_iacq_data & io_inner_acquire_valid;
  assign T230 = T59 & T231;
  assign T231 = T232[1'h0:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = 2'h0;
  assign T234 = T238 ? io_inner_acquire_bits_data : T235;
  assign T235 = T236 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T236 = T229 & T237;
  assign T237 = T227[1'h1:1'h1];
  assign T238 = T59 & T239;
  assign T239 = T232[1'h1:1'h1];
  assign T240 = T241[1'h0:1'h0];
  assign T241 = oacq_data_cnt;
  assign oacq_data_cnt = T111 ? R107 : 2'h0;
  assign T242 = T255 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T243 = T247 ? io_inner_acquire_bits_data : T244;
  assign T244 = T245 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T245 = T229 & T246;
  assign T246 = T227[2'h2:2'h2];
  assign T247 = T59 & T248;
  assign T248 = T232[2'h2:2'h2];
  assign T249 = T253 ? io_inner_acquire_bits_data : T250;
  assign T250 = T251 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T251 = T229 & T252;
  assign T252 = T227[2'h3:2'h3];
  assign T253 = T59 & T254;
  assign T254 = T232[2'h3:2'h3];
  assign T255 = T241[1'h0:1'h0];
  assign T256 = T241[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T257 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T258 = state == 3'h1;
  assign io_outer_acquire_bits_union = T259;
  assign T259 = T258 ? oacq_probe_union : T260;
  assign T260 = T257 ? T267 : T261;
  assign T261 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T419;
  assign T419 = {4'h0, T262};
  assign T262 = {T263, 6'h0};
  assign T263 = {T266, T264};
  assign T264 = xact_union[4'h8:3'h6];
  assign T265 = T59 ? io_inner_acquire_bits_union : xact_union;
  assign T266 = xact_union[4'hc:4'h9];
  assign T267 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T268;
  assign T268 = {T269, 1'h1};
  assign T269 = 16'hffff;
  assign oacq_write_beat_union = T270;
  assign T270 = {T271, 1'h1};
  assign T271 = T288 ? T279 : T272;
  assign T272 = T274 ? T273 : 16'h0;
  assign T273 = xact_union[5'h10:1'h1];
  assign T274 = T277 | T275;
  assign T275 = xact_is_builtin_type & T276;
  assign T276 = xact_a_type == 3'h2;
  assign T277 = xact_is_builtin_type & T278;
  assign T278 = xact_a_type == 3'h3;
  assign T279 = T280;
  assign T280 = {T286, T281};
  assign T281 = 8'h0 - T420;
  assign T420 = {7'h0, T282};
  assign T282 = T283[1'h0:1'h0];
  assign T283 = 1'h1 << T284;
  assign T284 = T285[2'h3:2'h3];
  assign T285 = xact_union[4'hc:4'h9];
  assign T286 = 8'h0 - T421;
  assign T421 = {7'h0, T287};
  assign T287 = T283[1'h1:1'h1];
  assign T288 = xact_is_builtin_type & T289;
  assign T289 = xact_a_type == 3'h4;
  assign oacq_probe_union = T290;
  assign T290 = {T291, 1'h1};
  assign T291 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T292;
  assign T292 = T258 ? oacq_probe_a_type : T293;
  assign T293 = T257 ? T295 : T294;
  assign T294 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T295 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T296;
  assign T296 = T258 ? oacq_probe_is_builtin_type : T297;
  assign T297 = T257 ? T299 : T298;
  assign T298 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T299 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T300;
  assign T300 = T258 ? oacq_probe_addr_beat : T301;
  assign T301 = T257 ? T304 : T302;
  assign T302 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T303 = T59 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T304 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T305;
  assign T305 = T258 ? oacq_probe_client_xact_id : T306;
  assign T306 = T257 ? T308 : T307;
  assign T307 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h3;
  assign oacq_read_beat_client_xact_id = 4'h3;
  assign T308 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h3;
  assign oacq_write_beat_client_xact_id = 4'h3;
  assign oacq_probe_client_xact_id = 4'h3;
  assign io_outer_acquire_bits_addr_block = T309;
  assign T309 = T258 ? oacq_probe_addr_block : T310;
  assign T310 = T257 ? T312 : T311;
  assign T311 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T312 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T313;
  assign T313 = T124 ? T340 : T314;
  assign T314 = T121 ? T315 : T114;
  assign T315 = T339 & T316;
  assign T316 = T338 | T317;
  assign T317 = T322 & T318;
  assign T318 = T319 - 1'h1;
  assign T319 = 1'h1 << T320;
  assign T320 = T321 + 2'h1;
  assign T321 = oacq_data_cnt - oacq_data_cnt;
  assign T322 = iacq_data_valid >> oacq_data_cnt;
  assign T422 = reset ? 4'h0 : T323;
  assign T323 = T59 ? T331 : T324;
  assign T324 = T229 ? T325 : iacq_data_valid;
  assign T325 = T329 | T326;
  assign T326 = T423 & T327;
  assign T327 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T423 = T328 ? 4'hf : 4'h0;
  assign T328 = 1'h1;
  assign T329 = iacq_data_valid & T330;
  assign T330 = ~ T327;
  assign T331 = T332 << io_inner_acquire_bits_addr_beat;
  assign T332 = io_inner_acquire_bits_is_builtin_type & T333;
  assign T333 = T335 | T334;
  assign T334 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T335 = T337 | T336;
  assign T336 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T337 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T338 = collect_iacq_data ^ 1'h1;
  assign T339 = pending_ognt_ack ^ 1'h1;
  assign T340 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T341;
  assign T341 = T102 ? T342 : 1'h0;
  assign T342 = T343 | io_outer_acquire_ready;
  assign T343 = T344 ^ 1'h1;
  assign T344 = T346 | T345;
  assign T345 = 3'h2 == io_inner_release_bits_r_type;
  assign T346 = T348 | T347;
  assign T347 = 3'h1 == io_inner_release_bits_r_type;
  assign T348 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T349;
  assign T349 = T424;
  assign T424 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T356;
  assign T356 = T357;
  assign T357 = xact_is_builtin_type ? T362 : T358;
  assign T358 = T361 ? 2'h1 : T359;
  assign T359 = T360 ? 2'h0 : 2'h2;
  assign T360 = xact_a_type == 3'h1;
  assign T361 = xact_a_type == 3'h0;
  assign T362 = T371 ? 2'h2 : T363;
  assign T363 = T370 ? 2'h0 : T364;
  assign T364 = T369 ? 2'h2 : T365;
  assign T365 = T368 ? 2'h0 : T366;
  assign T366 = T367 ? 2'h0 : 2'h2;
  assign T367 = xact_a_type == 3'h4;
  assign T368 = xact_a_type == 3'h2;
  assign T369 = xact_a_type == 3'h0;
  assign T370 = xact_a_type == 3'h3;
  assign T371 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T372;
  assign T372 = xact_addr_block;
  assign io_inner_probe_valid = T373;
  assign T373 = T102 ? T374 : 1'h0;
  assign T374 = pending_probes != 1'h0;
  assign T425 = T426[1'h0:1'h0];
  assign T426 = reset ? 4'h0 : T350;
  assign T350 = T355 ? T428 : T351;
  assign T351 = T91 ? mask_incoherent : T427;
  assign T427 = {3'h0, pending_probes};
  assign T428 = {2'h0, T352};
  assign T352 = T429 & T353;
  assign T353 = ~ T354;
  assign T354 = 1'h1 << 1'h0;
  assign T429 = {1'h0, pending_probes};
  assign T355 = T102 & io_inner_probe_ready;
  assign io_inner_finish_ready = T150;
  assign io_inner_grant_bits_client_id = T375;
  assign T375 = xact_client_id;
  assign io_inner_grant_bits_data = T376;
  assign T376 = 4'h0;
  assign io_inner_grant_bits_g_type = T377;
  assign T377 = T430;
  assign T430 = {1'h0, T378};
  assign T378 = xact_is_builtin_type ? T381 : T431;
  assign T431 = {1'h0, T379};
  assign T379 = T380 ? 2'h0 : 2'h1;
  assign T380 = xact_a_type == 3'h0;
  assign T381 = T392 ? 3'h4 : T382;
  assign T382 = T391 ? 3'h5 : T383;
  assign T383 = T390 ? 3'h3 : T384;
  assign T384 = T389 ? 3'h3 : T385;
  assign T385 = T388 ? 3'h4 : T386;
  assign T386 = T387 ? 3'h1 : 3'h3;
  assign T387 = xact_a_type == 3'h5;
  assign T388 = xact_a_type == 3'h4;
  assign T389 = xact_a_type == 3'h3;
  assign T390 = xact_a_type == 3'h2;
  assign T391 = xact_a_type == 3'h1;
  assign T392 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T393;
  assign T393 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T394;
  assign T394 = 4'h3;
  assign io_inner_grant_bits_client_xact_id = T395;
  assign T395 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T396;
  assign T396 = 2'h0;
  assign io_inner_grant_valid = T397;
  assign T397 = T148 ? 1'h1 : T398;
  assign T398 = T142 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T399;
  assign T399 = T60 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T185 <= 1'b1;
  if(!T186 && T185 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T175 <= 1'b1;
  if(!T176 && T175 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T151 <= 1'b1;
  if(!T152 && T151 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= 3'h0;
    end else if(T147) begin
      state <= T143;
    end else if(T129) begin
      state <= T125;
    end else if(T122) begin
      state <= 3'h5;
    end else if(T120) begin
      state <= T119;
    end else if(T117) begin
      state <= T115;
    end else if(T76) begin
      state <= T61;
    end else if(T59) begin
      state <= T19;
    end
    if(T59) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T59) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T406;
    if(reset) begin
      R107 <= 2'h0;
    end else if(T110) begin
      R107 <= T109;
    end
    if(reset) begin
      R133 <= 2'h0;
    end else if(T136) begin
      R133 <= T135;
    end
    if(T59) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T59) begin
      collect_iacq_data <= T172;
    end else if(T162) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R166 <= 2'h0;
    end else if(T169) begin
      R166 <= T168;
    end
    if(T59) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T59) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T120) begin
      pending_ognt_ack <= 1'h1;
    end else if(T103) begin
      pending_ognt_ack <= 1'h1;
    end else if(T211) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T230) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T225) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T238) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T236) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T247) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T245) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T253) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T251) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T59) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T59) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T59) begin
      iacq_data_valid <= T331;
    end else if(T229) begin
      iacq_data_valid <= T325;
    end
    pending_probes <= T425;
  end
endmodule

module BroadcastAcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T400;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T401;
  wire[2:0] T25;
  wire[2:0] T402;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire pending_outer_write_;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[3:0] mask_incoherent;
  wire[3:0] T403;
  wire T51;
  wire T52;
  wire[3:0] mask_self;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T404;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T405;
  wire T58;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[2:0] T62;
  wire pending_outer_read;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire pending_outer_write;
  wire T69;
  wire T70;
  reg [2:0] xact_a_type;
  wire[2:0] T71;
  wire T72;
  wire T73;
  wire T74;
  reg  xact_is_builtin_type;
  wire T75;
  wire T76;
  wire T77;
  reg  release_count;
  wire T406;
  wire[2:0] T407;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T408;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire T85;
  wire[1:0] T409;
  wire T86;
  wire[2:0] T410;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T411;
  wire T90;
  wire T91;
  wire[2:0] T412;
  wire T92;
  wire[2:0] T413;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire oacq_data_done;
  wire T104;
  wire T105;
  wire T106;
  reg [1:0] R107;
  wire[1:0] T414;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire[2:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire ignt_data_done;
  wire T130;
  wire T131;
  wire T132;
  reg [1:0] R133;
  wire[1:0] T415;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire[2:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  reg[0:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire T159;
  reg  collect_iacq_data;
  wire T416;
  wire T160;
  wire T161;
  wire T162;
  wire iacq_data_done;
  wire T163;
  wire T164;
  wire T165;
  reg [1:0] R166;
  wire[1:0] T417;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  reg[0:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  reg [1:0] xact_client_id;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  reg[0:0] T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  reg [25:0] xact_addr_block;
  wire[25:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  reg  pending_ognt_ack;
  wire T418;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[3:0] T214;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[3:0] T220;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T221;
  wire[3:0] T222;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T223;
  wire[3:0] T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[1:0] T228;
  wire T229;
  wire T230;
  wire T231;
  wire[3:0] T232;
  wire[1:0] T233;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T234;
  wire[3:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[1:0] T241;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T242;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T243;
  wire[3:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T249;
  wire[3:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] oacq_write_beat_data;
  wire T257;
  wire[3:0] oacq_probe_data;
  wire T258;
  wire[16:0] T259;
  wire[16:0] T260;
  wire[16:0] T261;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T419;
  wire[12:0] T262;
  wire[6:0] T263;
  wire[2:0] T264;
  reg [16:0] xact_union;
  wire[16:0] T265;
  wire[3:0] T266;
  wire[16:0] T267;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T268;
  wire[15:0] T269;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T270;
  wire[15:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[15:0] T279;
  wire[15:0] T280;
  wire[7:0] T281;
  wire[7:0] T420;
  wire T282;
  wire[1:0] T283;
  wire T284;
  wire[3:0] T285;
  wire[7:0] T286;
  wire[7:0] T421;
  wire T287;
  wire T288;
  wire T289;
  wire[16:0] oacq_probe_union;
  wire[16:0] T290;
  wire[15:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[2:0] T294;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T295;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T296;
  wire T297;
  wire T298;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T299;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T303;
  wire[1:0] T304;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T308;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T309;
  wire[25:0] T310;
  wire[25:0] T311;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T312;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire[1:0] T321;
  wire T322;
  reg [3:0] iacq_data_valid;
  wire[3:0] T422;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[3:0] T326;
  wire[3:0] T327;
  wire[3:0] T423;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire[1:0] T349;
  wire[1:0] T424;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[1:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[25:0] T372;
  wire T373;
  wire T374;
  reg  pending_probes;
  wire T425;
  wire[3:0] T426;
  wire[3:0] T350;
  wire[3:0] T351;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[1:0] T352;
  wire T353;
  wire T354;
  wire[1:0] T429;
  wire T355;
  wire[1:0] T375;
  wire[3:0] T376;
  wire[3:0] T377;
  wire[3:0] T430;
  wire[2:0] T378;
  wire[2:0] T431;
  wire[1:0] T379;
  wire T380;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] T384;
  wire[2:0] T385;
  wire[2:0] T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[3:0] T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire T397;
  wire T398;
  wire T399;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R107 = {1{$random}};
    R133 = {1{$random}};
    T151 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R166 = {1{$random}};
    T175 = 1'b0;
    xact_client_id = {1{$random}};
    T185 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T400 = reset ? 3'h0 : T11;
  assign T11 = T149 ? 3'h0 : T12;
  assign T12 = T147 ? T143 : T13;
  assign T13 = T129 ? T125 : T14;
  assign T14 = T122 ? 3'h5 : T15;
  assign T15 = T120 ? T119 : T16;
  assign T16 = T117 ? T115 : T17;
  assign T17 = T76 ? T61 : T18;
  assign T18 = T59 ? T19 : state;
  assign T19 = T50 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T44 ? T41 : T22;
  assign T22 = T40 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T401;
  assign T401 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T402;
  assign T402 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T39 ? 3'h4 : T29;
  assign T29 = T38 ? 3'h5 : T30;
  assign T30 = T37 ? 3'h3 : T31;
  assign T31 = T36 ? 3'h3 : T32;
  assign T32 = T35 ? 3'h4 : T33;
  assign T33 = T34 ? 3'h1 : 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h5;
  assign T35 = io_inner_acquire_bits_a_type == 3'h4;
  assign T36 = io_inner_acquire_bits_a_type == 3'h3;
  assign T37 = io_inner_acquire_bits_a_type == 3'h2;
  assign T38 = io_inner_acquire_bits_a_type == 3'h1;
  assign T39 = io_inner_acquire_bits_a_type == 3'h0;
  assign T40 = 4'h0 == T24;
  assign T41 = T43 | T42;
  assign T42 = 4'h4 == T24;
  assign T43 = 4'h5 == T24;
  assign T44 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T45;
  assign T45 = T47 | T46;
  assign T46 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T49 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T50 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T403;
  assign T403 = {3'h0, T51};
  assign T51 = ~ T52;
  assign T52 = io_incoherent_0;
  assign mask_self = T56 | T53;
  assign T53 = T404 & T54;
  assign T54 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T404 = T55 ? 4'hf : 4'h0;
  assign T55 = 1'h0;
  assign T56 = T405 & T57;
  assign T57 = ~ T54;
  assign T405 = {3'h0, T58};
  assign T58 = 1'h1;
  assign T59 = T60 & io_inner_acquire_valid;
  assign T60 = 3'h0 == state;
  assign T61 = pending_outer_write ? 3'h3 : T62;
  assign T62 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T66 : T63;
  assign T63 = T65 | T64;
  assign T64 = 4'h1 == io_inner_grant_bits_g_type;
  assign T65 = 4'h0 == io_inner_grant_bits_g_type;
  assign T66 = T68 | T67;
  assign T67 = 4'h4 == io_inner_grant_bits_g_type;
  assign T68 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T69;
  assign T69 = T72 | T70;
  assign T70 = 3'h4 == xact_a_type;
  assign T71 = T59 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T72 = T74 | T73;
  assign T73 = 3'h3 == xact_a_type;
  assign T74 = 3'h2 == xact_a_type;
  assign T75 = T59 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T76 = T103 & T77;
  assign T77 = release_count == 1'h1;
  assign T406 = T407[1'h0:1'h0];
  assign T407 = reset ? 3'h0 : T78;
  assign T78 = T94 ? T413 : T79;
  assign T79 = T103 ? T412 : T80;
  assign T80 = T91 ? T81 : T408;
  assign T408 = {2'h0, release_count};
  assign T81 = T410 + T82;
  assign T82 = {1'h0, T83};
  assign T83 = T409 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = mask_incoherent[2'h3:2'h3];
  assign T409 = {1'h0, T86};
  assign T86 = mask_incoherent[2'h2:2'h2];
  assign T410 = {1'h0, T87};
  assign T87 = T411 + T88;
  assign T88 = {1'h0, T89};
  assign T89 = mask_incoherent[1'h1:1'h1];
  assign T411 = {1'h0, T90};
  assign T90 = mask_incoherent[1'h0:1'h0];
  assign T91 = T59 & T50;
  assign T412 = {2'h0, T92};
  assign T92 = release_count - 1'h1;
  assign T413 = {2'h0, T93};
  assign T93 = release_count - 1'h1;
  assign T94 = T101 & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = T98 | T97;
  assign T97 = 3'h2 == io_inner_release_bits_r_type;
  assign T98 = T100 | T99;
  assign T99 = 3'h1 == io_inner_release_bits_r_type;
  assign T100 = 3'h0 == io_inner_release_bits_r_type;
  assign T101 = T102 & io_inner_release_valid;
  assign T102 = 3'h1 == state;
  assign T103 = T113 & oacq_data_done;
  assign oacq_data_done = T111 ? T105 : T104;
  assign T104 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T105 = T110 & T106;
  assign T106 = R107 == 2'h3;
  assign T414 = reset ? 2'h0 : T108;
  assign T108 = T110 ? T109 : R107;
  assign T109 = R107 + 2'h1;
  assign T110 = T104 & T111;
  assign T111 = io_outer_acquire_bits_is_builtin_type & T112;
  assign T112 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T113 = T114 & io_outer_acquire_ready;
  assign T114 = T101 & T96;
  assign T115 = pending_outer_write ? 3'h3 : T116;
  assign T116 = pending_outer_read ? 3'h2 : 3'h4;
  assign T117 = T94 & T118;
  assign T118 = release_count == 1'h1;
  assign T119 = pending_outer_read ? 3'h2 : 3'h5;
  assign T120 = T121 & oacq_data_done;
  assign T121 = 3'h3 == state;
  assign T122 = T124 & T123;
  assign T123 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T124 = 3'h2 == state;
  assign T125 = T126 ? 3'h6 : 3'h0;
  assign T126 = T127 ^ 1'h1;
  assign T127 = io_inner_grant_bits_is_builtin_type & T128;
  assign T128 = io_inner_grant_bits_g_type == 4'h0;
  assign T129 = T142 & ignt_data_done;
  assign ignt_data_done = T137 ? T131 : T130;
  assign T130 = io_inner_grant_ready & io_inner_grant_valid;
  assign T131 = T136 & T132;
  assign T132 = R133 == 2'h3;
  assign T415 = reset ? 2'h0 : T134;
  assign T134 = T136 ? T135 : R133;
  assign T135 = R133 + 2'h1;
  assign T136 = T130 & T137;
  assign T137 = io_inner_grant_bits_is_builtin_type ? T141 : T138;
  assign T138 = T140 | T139;
  assign T139 = 4'h1 == io_inner_grant_bits_g_type;
  assign T140 = 4'h0 == io_inner_grant_bits_g_type;
  assign T141 = 4'h5 == io_inner_grant_bits_g_type;
  assign T142 = 3'h5 == state;
  assign T143 = T144 ? 3'h6 : 3'h0;
  assign T144 = T145 ^ 1'h1;
  assign T145 = io_inner_grant_bits_is_builtin_type & T146;
  assign T146 = io_inner_grant_bits_g_type == 4'h0;
  assign T147 = T148 & io_inner_grant_ready;
  assign T148 = 3'h4 == state;
  assign T149 = T150 & io_inner_finish_valid;
  assign T150 = 3'h6 == state;
  assign T152 = T153 | reset;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T157 & T155;
  assign T155 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T156 = T59 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T157 = T159 & T158;
  assign T158 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T159 = T174 & collect_iacq_data;
  assign T416 = reset ? 1'h0 : T160;
  assign T160 = T59 ? T172 : T161;
  assign T161 = T162 ? 1'h0 : collect_iacq_data;
  assign T162 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T170 ? T164 : T163;
  assign T163 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T164 = T169 & T165;
  assign T165 = R166 == 2'h3;
  assign T417 = reset ? 2'h0 : T167;
  assign T167 = T169 ? T168 : R166;
  assign T168 = R166 + 2'h1;
  assign T169 = T163 & T170;
  assign T170 = io_inner_acquire_bits_is_builtin_type & T171;
  assign T171 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = state != 3'h0;
  assign T176 = T177 | reset;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T181 & T179;
  assign T179 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T180 = T59 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T181 = T183 & T182;
  assign T182 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T183 = T184 & collect_iacq_data;
  assign T184 = state != 3'h0;
  assign T186 = T187 | reset;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T192 & T189;
  assign T189 = T191 | T190;
  assign T190 = 3'h5 == xact_a_type;
  assign T191 = 3'h4 == xact_a_type;
  assign T192 = T193 & xact_is_builtin_type;
  assign T193 = state != 3'h0;
  assign io_has_release_match = T194;
  assign T194 = T196 & T195;
  assign T195 = state == 3'h1;
  assign T196 = T198 & T197;
  assign T197 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T198 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T199 = T59 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T200;
  assign T200 = T201 & collect_iacq_data;
  assign T201 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T202;
  assign T202 = T204 & T203;
  assign T203 = collect_iacq_data ^ 1'h1;
  assign T204 = T206 & T205;
  assign T205 = state != 3'h0;
  assign T206 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T207;
  assign T207 = T142 ? io_inner_grant_ready : pending_ognt_ack;
  assign T418 = reset ? 1'h0 : T208;
  assign T208 = T120 ? 1'h1 : T209;
  assign T209 = T103 ? 1'h1 : T210;
  assign T210 = T211 ? 1'h0 : pending_ognt_ack;
  assign T211 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T212;
  assign T212 = T258 ? oacq_probe_data : T213;
  assign T213 = T257 ? T220 : T214;
  assign T214 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T215;
  assign T215 = T217 | T216;
  assign T216 = 3'h4 == xact_a_type;
  assign T217 = T219 | T218;
  assign T218 = 3'h0 == xact_a_type;
  assign T219 = 3'h2 == xact_a_type;
  assign T220 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T221;
  assign T221 = T256 ? T242 : T222;
  assign T222 = T240 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T223 = T230 ? io_inner_acquire_bits_data : T224;
  assign T224 = T225 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T225 = T229 & T226;
  assign T226 = T227[1'h0:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = io_inner_acquire_bits_addr_beat;
  assign T229 = collect_iacq_data & io_inner_acquire_valid;
  assign T230 = T59 & T231;
  assign T231 = T232[1'h0:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = 2'h0;
  assign T234 = T238 ? io_inner_acquire_bits_data : T235;
  assign T235 = T236 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T236 = T229 & T237;
  assign T237 = T227[1'h1:1'h1];
  assign T238 = T59 & T239;
  assign T239 = T232[1'h1:1'h1];
  assign T240 = T241[1'h0:1'h0];
  assign T241 = oacq_data_cnt;
  assign oacq_data_cnt = T111 ? R107 : 2'h0;
  assign T242 = T255 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T243 = T247 ? io_inner_acquire_bits_data : T244;
  assign T244 = T245 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T245 = T229 & T246;
  assign T246 = T227[2'h2:2'h2];
  assign T247 = T59 & T248;
  assign T248 = T232[2'h2:2'h2];
  assign T249 = T253 ? io_inner_acquire_bits_data : T250;
  assign T250 = T251 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T251 = T229 & T252;
  assign T252 = T227[2'h3:2'h3];
  assign T253 = T59 & T254;
  assign T254 = T232[2'h3:2'h3];
  assign T255 = T241[1'h0:1'h0];
  assign T256 = T241[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T257 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T258 = state == 3'h1;
  assign io_outer_acquire_bits_union = T259;
  assign T259 = T258 ? oacq_probe_union : T260;
  assign T260 = T257 ? T267 : T261;
  assign T261 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T419;
  assign T419 = {4'h0, T262};
  assign T262 = {T263, 6'h0};
  assign T263 = {T266, T264};
  assign T264 = xact_union[4'h8:3'h6];
  assign T265 = T59 ? io_inner_acquire_bits_union : xact_union;
  assign T266 = xact_union[4'hc:4'h9];
  assign T267 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T268;
  assign T268 = {T269, 1'h1};
  assign T269 = 16'hffff;
  assign oacq_write_beat_union = T270;
  assign T270 = {T271, 1'h1};
  assign T271 = T288 ? T279 : T272;
  assign T272 = T274 ? T273 : 16'h0;
  assign T273 = xact_union[5'h10:1'h1];
  assign T274 = T277 | T275;
  assign T275 = xact_is_builtin_type & T276;
  assign T276 = xact_a_type == 3'h2;
  assign T277 = xact_is_builtin_type & T278;
  assign T278 = xact_a_type == 3'h3;
  assign T279 = T280;
  assign T280 = {T286, T281};
  assign T281 = 8'h0 - T420;
  assign T420 = {7'h0, T282};
  assign T282 = T283[1'h0:1'h0];
  assign T283 = 1'h1 << T284;
  assign T284 = T285[2'h3:2'h3];
  assign T285 = xact_union[4'hc:4'h9];
  assign T286 = 8'h0 - T421;
  assign T421 = {7'h0, T287};
  assign T287 = T283[1'h1:1'h1];
  assign T288 = xact_is_builtin_type & T289;
  assign T289 = xact_a_type == 3'h4;
  assign oacq_probe_union = T290;
  assign T290 = {T291, 1'h1};
  assign T291 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T292;
  assign T292 = T258 ? oacq_probe_a_type : T293;
  assign T293 = T257 ? T295 : T294;
  assign T294 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T295 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T296;
  assign T296 = T258 ? oacq_probe_is_builtin_type : T297;
  assign T297 = T257 ? T299 : T298;
  assign T298 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T299 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T300;
  assign T300 = T258 ? oacq_probe_addr_beat : T301;
  assign T301 = T257 ? T304 : T302;
  assign T302 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T303 = T59 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T304 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T305;
  assign T305 = T258 ? oacq_probe_client_xact_id : T306;
  assign T306 = T257 ? T308 : T307;
  assign T307 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h4;
  assign oacq_read_beat_client_xact_id = 4'h4;
  assign T308 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h4;
  assign oacq_write_beat_client_xact_id = 4'h4;
  assign oacq_probe_client_xact_id = 4'h4;
  assign io_outer_acquire_bits_addr_block = T309;
  assign T309 = T258 ? oacq_probe_addr_block : T310;
  assign T310 = T257 ? T312 : T311;
  assign T311 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T312 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T313;
  assign T313 = T124 ? T340 : T314;
  assign T314 = T121 ? T315 : T114;
  assign T315 = T339 & T316;
  assign T316 = T338 | T317;
  assign T317 = T322 & T318;
  assign T318 = T319 - 1'h1;
  assign T319 = 1'h1 << T320;
  assign T320 = T321 + 2'h1;
  assign T321 = oacq_data_cnt - oacq_data_cnt;
  assign T322 = iacq_data_valid >> oacq_data_cnt;
  assign T422 = reset ? 4'h0 : T323;
  assign T323 = T59 ? T331 : T324;
  assign T324 = T229 ? T325 : iacq_data_valid;
  assign T325 = T329 | T326;
  assign T326 = T423 & T327;
  assign T327 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T423 = T328 ? 4'hf : 4'h0;
  assign T328 = 1'h1;
  assign T329 = iacq_data_valid & T330;
  assign T330 = ~ T327;
  assign T331 = T332 << io_inner_acquire_bits_addr_beat;
  assign T332 = io_inner_acquire_bits_is_builtin_type & T333;
  assign T333 = T335 | T334;
  assign T334 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T335 = T337 | T336;
  assign T336 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T337 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T338 = collect_iacq_data ^ 1'h1;
  assign T339 = pending_ognt_ack ^ 1'h1;
  assign T340 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T341;
  assign T341 = T102 ? T342 : 1'h0;
  assign T342 = T343 | io_outer_acquire_ready;
  assign T343 = T344 ^ 1'h1;
  assign T344 = T346 | T345;
  assign T345 = 3'h2 == io_inner_release_bits_r_type;
  assign T346 = T348 | T347;
  assign T347 = 3'h1 == io_inner_release_bits_r_type;
  assign T348 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T349;
  assign T349 = T424;
  assign T424 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T356;
  assign T356 = T357;
  assign T357 = xact_is_builtin_type ? T362 : T358;
  assign T358 = T361 ? 2'h1 : T359;
  assign T359 = T360 ? 2'h0 : 2'h2;
  assign T360 = xact_a_type == 3'h1;
  assign T361 = xact_a_type == 3'h0;
  assign T362 = T371 ? 2'h2 : T363;
  assign T363 = T370 ? 2'h0 : T364;
  assign T364 = T369 ? 2'h2 : T365;
  assign T365 = T368 ? 2'h0 : T366;
  assign T366 = T367 ? 2'h0 : 2'h2;
  assign T367 = xact_a_type == 3'h4;
  assign T368 = xact_a_type == 3'h2;
  assign T369 = xact_a_type == 3'h0;
  assign T370 = xact_a_type == 3'h3;
  assign T371 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T372;
  assign T372 = xact_addr_block;
  assign io_inner_probe_valid = T373;
  assign T373 = T102 ? T374 : 1'h0;
  assign T374 = pending_probes != 1'h0;
  assign T425 = T426[1'h0:1'h0];
  assign T426 = reset ? 4'h0 : T350;
  assign T350 = T355 ? T428 : T351;
  assign T351 = T91 ? mask_incoherent : T427;
  assign T427 = {3'h0, pending_probes};
  assign T428 = {2'h0, T352};
  assign T352 = T429 & T353;
  assign T353 = ~ T354;
  assign T354 = 1'h1 << 1'h0;
  assign T429 = {1'h0, pending_probes};
  assign T355 = T102 & io_inner_probe_ready;
  assign io_inner_finish_ready = T150;
  assign io_inner_grant_bits_client_id = T375;
  assign T375 = xact_client_id;
  assign io_inner_grant_bits_data = T376;
  assign T376 = 4'h0;
  assign io_inner_grant_bits_g_type = T377;
  assign T377 = T430;
  assign T430 = {1'h0, T378};
  assign T378 = xact_is_builtin_type ? T381 : T431;
  assign T431 = {1'h0, T379};
  assign T379 = T380 ? 2'h0 : 2'h1;
  assign T380 = xact_a_type == 3'h0;
  assign T381 = T392 ? 3'h4 : T382;
  assign T382 = T391 ? 3'h5 : T383;
  assign T383 = T390 ? 3'h3 : T384;
  assign T384 = T389 ? 3'h3 : T385;
  assign T385 = T388 ? 3'h4 : T386;
  assign T386 = T387 ? 3'h1 : 3'h3;
  assign T387 = xact_a_type == 3'h5;
  assign T388 = xact_a_type == 3'h4;
  assign T389 = xact_a_type == 3'h3;
  assign T390 = xact_a_type == 3'h2;
  assign T391 = xact_a_type == 3'h1;
  assign T392 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T393;
  assign T393 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T394;
  assign T394 = 4'h4;
  assign io_inner_grant_bits_client_xact_id = T395;
  assign T395 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T396;
  assign T396 = 2'h0;
  assign io_inner_grant_valid = T397;
  assign T397 = T148 ? 1'h1 : T398;
  assign T398 = T142 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T399;
  assign T399 = T60 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T185 <= 1'b1;
  if(!T186 && T185 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T175 <= 1'b1;
  if(!T176 && T175 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T151 <= 1'b1;
  if(!T152 && T151 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= 3'h0;
    end else if(T147) begin
      state <= T143;
    end else if(T129) begin
      state <= T125;
    end else if(T122) begin
      state <= 3'h5;
    end else if(T120) begin
      state <= T119;
    end else if(T117) begin
      state <= T115;
    end else if(T76) begin
      state <= T61;
    end else if(T59) begin
      state <= T19;
    end
    if(T59) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T59) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T406;
    if(reset) begin
      R107 <= 2'h0;
    end else if(T110) begin
      R107 <= T109;
    end
    if(reset) begin
      R133 <= 2'h0;
    end else if(T136) begin
      R133 <= T135;
    end
    if(T59) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T59) begin
      collect_iacq_data <= T172;
    end else if(T162) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R166 <= 2'h0;
    end else if(T169) begin
      R166 <= T168;
    end
    if(T59) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T59) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T120) begin
      pending_ognt_ack <= 1'h1;
    end else if(T103) begin
      pending_ognt_ack <= 1'h1;
    end else if(T211) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T230) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T225) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T238) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T236) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T247) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T245) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T253) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T251) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T59) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T59) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T59) begin
      iacq_data_valid <= T331;
    end else if(T229) begin
      iacq_data_valid <= T325;
    end
    pending_probes <= T425;
  end
endmodule

module BroadcastAcquireTracker_4(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T400;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T401;
  wire[2:0] T25;
  wire[2:0] T402;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire pending_outer_write_;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[3:0] mask_incoherent;
  wire[3:0] T403;
  wire T51;
  wire T52;
  wire[3:0] mask_self;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T404;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T405;
  wire T58;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[2:0] T62;
  wire pending_outer_read;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire pending_outer_write;
  wire T69;
  wire T70;
  reg [2:0] xact_a_type;
  wire[2:0] T71;
  wire T72;
  wire T73;
  wire T74;
  reg  xact_is_builtin_type;
  wire T75;
  wire T76;
  wire T77;
  reg  release_count;
  wire T406;
  wire[2:0] T407;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T408;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire T85;
  wire[1:0] T409;
  wire T86;
  wire[2:0] T410;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T411;
  wire T90;
  wire T91;
  wire[2:0] T412;
  wire T92;
  wire[2:0] T413;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire oacq_data_done;
  wire T104;
  wire T105;
  wire T106;
  reg [1:0] R107;
  wire[1:0] T414;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire[2:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire ignt_data_done;
  wire T130;
  wire T131;
  wire T132;
  reg [1:0] R133;
  wire[1:0] T415;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire[2:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  reg[0:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire T159;
  reg  collect_iacq_data;
  wire T416;
  wire T160;
  wire T161;
  wire T162;
  wire iacq_data_done;
  wire T163;
  wire T164;
  wire T165;
  reg [1:0] R166;
  wire[1:0] T417;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  reg[0:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  reg [1:0] xact_client_id;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  reg[0:0] T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  reg [25:0] xact_addr_block;
  wire[25:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  reg  pending_ognt_ack;
  wire T418;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[3:0] T214;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[3:0] T220;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T221;
  wire[3:0] T222;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T223;
  wire[3:0] T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[1:0] T228;
  wire T229;
  wire T230;
  wire T231;
  wire[3:0] T232;
  wire[1:0] T233;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T234;
  wire[3:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[1:0] T241;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T242;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T243;
  wire[3:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T249;
  wire[3:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] oacq_write_beat_data;
  wire T257;
  wire[3:0] oacq_probe_data;
  wire T258;
  wire[16:0] T259;
  wire[16:0] T260;
  wire[16:0] T261;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T419;
  wire[12:0] T262;
  wire[6:0] T263;
  wire[2:0] T264;
  reg [16:0] xact_union;
  wire[16:0] T265;
  wire[3:0] T266;
  wire[16:0] T267;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T268;
  wire[15:0] T269;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T270;
  wire[15:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[15:0] T279;
  wire[15:0] T280;
  wire[7:0] T281;
  wire[7:0] T420;
  wire T282;
  wire[1:0] T283;
  wire T284;
  wire[3:0] T285;
  wire[7:0] T286;
  wire[7:0] T421;
  wire T287;
  wire T288;
  wire T289;
  wire[16:0] oacq_probe_union;
  wire[16:0] T290;
  wire[15:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[2:0] T294;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T295;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T296;
  wire T297;
  wire T298;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T299;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T303;
  wire[1:0] T304;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T308;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T309;
  wire[25:0] T310;
  wire[25:0] T311;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T312;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire[1:0] T321;
  wire T322;
  reg [3:0] iacq_data_valid;
  wire[3:0] T422;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[3:0] T326;
  wire[3:0] T327;
  wire[3:0] T423;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire[1:0] T349;
  wire[1:0] T424;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[1:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[25:0] T372;
  wire T373;
  wire T374;
  reg  pending_probes;
  wire T425;
  wire[3:0] T426;
  wire[3:0] T350;
  wire[3:0] T351;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[1:0] T352;
  wire T353;
  wire T354;
  wire[1:0] T429;
  wire T355;
  wire[1:0] T375;
  wire[3:0] T376;
  wire[3:0] T377;
  wire[3:0] T430;
  wire[2:0] T378;
  wire[2:0] T431;
  wire[1:0] T379;
  wire T380;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] T384;
  wire[2:0] T385;
  wire[2:0] T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[3:0] T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire T397;
  wire T398;
  wire T399;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R107 = {1{$random}};
    R133 = {1{$random}};
    T151 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R166 = {1{$random}};
    T175 = 1'b0;
    xact_client_id = {1{$random}};
    T185 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T400 = reset ? 3'h0 : T11;
  assign T11 = T149 ? 3'h0 : T12;
  assign T12 = T147 ? T143 : T13;
  assign T13 = T129 ? T125 : T14;
  assign T14 = T122 ? 3'h5 : T15;
  assign T15 = T120 ? T119 : T16;
  assign T16 = T117 ? T115 : T17;
  assign T17 = T76 ? T61 : T18;
  assign T18 = T59 ? T19 : state;
  assign T19 = T50 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T44 ? T41 : T22;
  assign T22 = T40 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T401;
  assign T401 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T402;
  assign T402 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T39 ? 3'h4 : T29;
  assign T29 = T38 ? 3'h5 : T30;
  assign T30 = T37 ? 3'h3 : T31;
  assign T31 = T36 ? 3'h3 : T32;
  assign T32 = T35 ? 3'h4 : T33;
  assign T33 = T34 ? 3'h1 : 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h5;
  assign T35 = io_inner_acquire_bits_a_type == 3'h4;
  assign T36 = io_inner_acquire_bits_a_type == 3'h3;
  assign T37 = io_inner_acquire_bits_a_type == 3'h2;
  assign T38 = io_inner_acquire_bits_a_type == 3'h1;
  assign T39 = io_inner_acquire_bits_a_type == 3'h0;
  assign T40 = 4'h0 == T24;
  assign T41 = T43 | T42;
  assign T42 = 4'h4 == T24;
  assign T43 = 4'h5 == T24;
  assign T44 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T45;
  assign T45 = T47 | T46;
  assign T46 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T49 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T50 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T403;
  assign T403 = {3'h0, T51};
  assign T51 = ~ T52;
  assign T52 = io_incoherent_0;
  assign mask_self = T56 | T53;
  assign T53 = T404 & T54;
  assign T54 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T404 = T55 ? 4'hf : 4'h0;
  assign T55 = 1'h0;
  assign T56 = T405 & T57;
  assign T57 = ~ T54;
  assign T405 = {3'h0, T58};
  assign T58 = 1'h1;
  assign T59 = T60 & io_inner_acquire_valid;
  assign T60 = 3'h0 == state;
  assign T61 = pending_outer_write ? 3'h3 : T62;
  assign T62 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T66 : T63;
  assign T63 = T65 | T64;
  assign T64 = 4'h1 == io_inner_grant_bits_g_type;
  assign T65 = 4'h0 == io_inner_grant_bits_g_type;
  assign T66 = T68 | T67;
  assign T67 = 4'h4 == io_inner_grant_bits_g_type;
  assign T68 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T69;
  assign T69 = T72 | T70;
  assign T70 = 3'h4 == xact_a_type;
  assign T71 = T59 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T72 = T74 | T73;
  assign T73 = 3'h3 == xact_a_type;
  assign T74 = 3'h2 == xact_a_type;
  assign T75 = T59 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T76 = T103 & T77;
  assign T77 = release_count == 1'h1;
  assign T406 = T407[1'h0:1'h0];
  assign T407 = reset ? 3'h0 : T78;
  assign T78 = T94 ? T413 : T79;
  assign T79 = T103 ? T412 : T80;
  assign T80 = T91 ? T81 : T408;
  assign T408 = {2'h0, release_count};
  assign T81 = T410 + T82;
  assign T82 = {1'h0, T83};
  assign T83 = T409 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = mask_incoherent[2'h3:2'h3];
  assign T409 = {1'h0, T86};
  assign T86 = mask_incoherent[2'h2:2'h2];
  assign T410 = {1'h0, T87};
  assign T87 = T411 + T88;
  assign T88 = {1'h0, T89};
  assign T89 = mask_incoherent[1'h1:1'h1];
  assign T411 = {1'h0, T90};
  assign T90 = mask_incoherent[1'h0:1'h0];
  assign T91 = T59 & T50;
  assign T412 = {2'h0, T92};
  assign T92 = release_count - 1'h1;
  assign T413 = {2'h0, T93};
  assign T93 = release_count - 1'h1;
  assign T94 = T101 & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = T98 | T97;
  assign T97 = 3'h2 == io_inner_release_bits_r_type;
  assign T98 = T100 | T99;
  assign T99 = 3'h1 == io_inner_release_bits_r_type;
  assign T100 = 3'h0 == io_inner_release_bits_r_type;
  assign T101 = T102 & io_inner_release_valid;
  assign T102 = 3'h1 == state;
  assign T103 = T113 & oacq_data_done;
  assign oacq_data_done = T111 ? T105 : T104;
  assign T104 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T105 = T110 & T106;
  assign T106 = R107 == 2'h3;
  assign T414 = reset ? 2'h0 : T108;
  assign T108 = T110 ? T109 : R107;
  assign T109 = R107 + 2'h1;
  assign T110 = T104 & T111;
  assign T111 = io_outer_acquire_bits_is_builtin_type & T112;
  assign T112 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T113 = T114 & io_outer_acquire_ready;
  assign T114 = T101 & T96;
  assign T115 = pending_outer_write ? 3'h3 : T116;
  assign T116 = pending_outer_read ? 3'h2 : 3'h4;
  assign T117 = T94 & T118;
  assign T118 = release_count == 1'h1;
  assign T119 = pending_outer_read ? 3'h2 : 3'h5;
  assign T120 = T121 & oacq_data_done;
  assign T121 = 3'h3 == state;
  assign T122 = T124 & T123;
  assign T123 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T124 = 3'h2 == state;
  assign T125 = T126 ? 3'h6 : 3'h0;
  assign T126 = T127 ^ 1'h1;
  assign T127 = io_inner_grant_bits_is_builtin_type & T128;
  assign T128 = io_inner_grant_bits_g_type == 4'h0;
  assign T129 = T142 & ignt_data_done;
  assign ignt_data_done = T137 ? T131 : T130;
  assign T130 = io_inner_grant_ready & io_inner_grant_valid;
  assign T131 = T136 & T132;
  assign T132 = R133 == 2'h3;
  assign T415 = reset ? 2'h0 : T134;
  assign T134 = T136 ? T135 : R133;
  assign T135 = R133 + 2'h1;
  assign T136 = T130 & T137;
  assign T137 = io_inner_grant_bits_is_builtin_type ? T141 : T138;
  assign T138 = T140 | T139;
  assign T139 = 4'h1 == io_inner_grant_bits_g_type;
  assign T140 = 4'h0 == io_inner_grant_bits_g_type;
  assign T141 = 4'h5 == io_inner_grant_bits_g_type;
  assign T142 = 3'h5 == state;
  assign T143 = T144 ? 3'h6 : 3'h0;
  assign T144 = T145 ^ 1'h1;
  assign T145 = io_inner_grant_bits_is_builtin_type & T146;
  assign T146 = io_inner_grant_bits_g_type == 4'h0;
  assign T147 = T148 & io_inner_grant_ready;
  assign T148 = 3'h4 == state;
  assign T149 = T150 & io_inner_finish_valid;
  assign T150 = 3'h6 == state;
  assign T152 = T153 | reset;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T157 & T155;
  assign T155 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T156 = T59 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T157 = T159 & T158;
  assign T158 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T159 = T174 & collect_iacq_data;
  assign T416 = reset ? 1'h0 : T160;
  assign T160 = T59 ? T172 : T161;
  assign T161 = T162 ? 1'h0 : collect_iacq_data;
  assign T162 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T170 ? T164 : T163;
  assign T163 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T164 = T169 & T165;
  assign T165 = R166 == 2'h3;
  assign T417 = reset ? 2'h0 : T167;
  assign T167 = T169 ? T168 : R166;
  assign T168 = R166 + 2'h1;
  assign T169 = T163 & T170;
  assign T170 = io_inner_acquire_bits_is_builtin_type & T171;
  assign T171 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = state != 3'h0;
  assign T176 = T177 | reset;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T181 & T179;
  assign T179 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T180 = T59 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T181 = T183 & T182;
  assign T182 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T183 = T184 & collect_iacq_data;
  assign T184 = state != 3'h0;
  assign T186 = T187 | reset;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T192 & T189;
  assign T189 = T191 | T190;
  assign T190 = 3'h5 == xact_a_type;
  assign T191 = 3'h4 == xact_a_type;
  assign T192 = T193 & xact_is_builtin_type;
  assign T193 = state != 3'h0;
  assign io_has_release_match = T194;
  assign T194 = T196 & T195;
  assign T195 = state == 3'h1;
  assign T196 = T198 & T197;
  assign T197 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T198 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T199 = T59 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T200;
  assign T200 = T201 & collect_iacq_data;
  assign T201 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T202;
  assign T202 = T204 & T203;
  assign T203 = collect_iacq_data ^ 1'h1;
  assign T204 = T206 & T205;
  assign T205 = state != 3'h0;
  assign T206 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T207;
  assign T207 = T142 ? io_inner_grant_ready : pending_ognt_ack;
  assign T418 = reset ? 1'h0 : T208;
  assign T208 = T120 ? 1'h1 : T209;
  assign T209 = T103 ? 1'h1 : T210;
  assign T210 = T211 ? 1'h0 : pending_ognt_ack;
  assign T211 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T212;
  assign T212 = T258 ? oacq_probe_data : T213;
  assign T213 = T257 ? T220 : T214;
  assign T214 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T215;
  assign T215 = T217 | T216;
  assign T216 = 3'h4 == xact_a_type;
  assign T217 = T219 | T218;
  assign T218 = 3'h0 == xact_a_type;
  assign T219 = 3'h2 == xact_a_type;
  assign T220 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T221;
  assign T221 = T256 ? T242 : T222;
  assign T222 = T240 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T223 = T230 ? io_inner_acquire_bits_data : T224;
  assign T224 = T225 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T225 = T229 & T226;
  assign T226 = T227[1'h0:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = io_inner_acquire_bits_addr_beat;
  assign T229 = collect_iacq_data & io_inner_acquire_valid;
  assign T230 = T59 & T231;
  assign T231 = T232[1'h0:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = 2'h0;
  assign T234 = T238 ? io_inner_acquire_bits_data : T235;
  assign T235 = T236 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T236 = T229 & T237;
  assign T237 = T227[1'h1:1'h1];
  assign T238 = T59 & T239;
  assign T239 = T232[1'h1:1'h1];
  assign T240 = T241[1'h0:1'h0];
  assign T241 = oacq_data_cnt;
  assign oacq_data_cnt = T111 ? R107 : 2'h0;
  assign T242 = T255 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T243 = T247 ? io_inner_acquire_bits_data : T244;
  assign T244 = T245 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T245 = T229 & T246;
  assign T246 = T227[2'h2:2'h2];
  assign T247 = T59 & T248;
  assign T248 = T232[2'h2:2'h2];
  assign T249 = T253 ? io_inner_acquire_bits_data : T250;
  assign T250 = T251 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T251 = T229 & T252;
  assign T252 = T227[2'h3:2'h3];
  assign T253 = T59 & T254;
  assign T254 = T232[2'h3:2'h3];
  assign T255 = T241[1'h0:1'h0];
  assign T256 = T241[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T257 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T258 = state == 3'h1;
  assign io_outer_acquire_bits_union = T259;
  assign T259 = T258 ? oacq_probe_union : T260;
  assign T260 = T257 ? T267 : T261;
  assign T261 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T419;
  assign T419 = {4'h0, T262};
  assign T262 = {T263, 6'h0};
  assign T263 = {T266, T264};
  assign T264 = xact_union[4'h8:3'h6];
  assign T265 = T59 ? io_inner_acquire_bits_union : xact_union;
  assign T266 = xact_union[4'hc:4'h9];
  assign T267 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T268;
  assign T268 = {T269, 1'h1};
  assign T269 = 16'hffff;
  assign oacq_write_beat_union = T270;
  assign T270 = {T271, 1'h1};
  assign T271 = T288 ? T279 : T272;
  assign T272 = T274 ? T273 : 16'h0;
  assign T273 = xact_union[5'h10:1'h1];
  assign T274 = T277 | T275;
  assign T275 = xact_is_builtin_type & T276;
  assign T276 = xact_a_type == 3'h2;
  assign T277 = xact_is_builtin_type & T278;
  assign T278 = xact_a_type == 3'h3;
  assign T279 = T280;
  assign T280 = {T286, T281};
  assign T281 = 8'h0 - T420;
  assign T420 = {7'h0, T282};
  assign T282 = T283[1'h0:1'h0];
  assign T283 = 1'h1 << T284;
  assign T284 = T285[2'h3:2'h3];
  assign T285 = xact_union[4'hc:4'h9];
  assign T286 = 8'h0 - T421;
  assign T421 = {7'h0, T287};
  assign T287 = T283[1'h1:1'h1];
  assign T288 = xact_is_builtin_type & T289;
  assign T289 = xact_a_type == 3'h4;
  assign oacq_probe_union = T290;
  assign T290 = {T291, 1'h1};
  assign T291 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T292;
  assign T292 = T258 ? oacq_probe_a_type : T293;
  assign T293 = T257 ? T295 : T294;
  assign T294 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T295 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T296;
  assign T296 = T258 ? oacq_probe_is_builtin_type : T297;
  assign T297 = T257 ? T299 : T298;
  assign T298 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T299 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T300;
  assign T300 = T258 ? oacq_probe_addr_beat : T301;
  assign T301 = T257 ? T304 : T302;
  assign T302 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T303 = T59 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T304 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T305;
  assign T305 = T258 ? oacq_probe_client_xact_id : T306;
  assign T306 = T257 ? T308 : T307;
  assign T307 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h5;
  assign oacq_read_beat_client_xact_id = 4'h5;
  assign T308 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h5;
  assign oacq_write_beat_client_xact_id = 4'h5;
  assign oacq_probe_client_xact_id = 4'h5;
  assign io_outer_acquire_bits_addr_block = T309;
  assign T309 = T258 ? oacq_probe_addr_block : T310;
  assign T310 = T257 ? T312 : T311;
  assign T311 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T312 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T313;
  assign T313 = T124 ? T340 : T314;
  assign T314 = T121 ? T315 : T114;
  assign T315 = T339 & T316;
  assign T316 = T338 | T317;
  assign T317 = T322 & T318;
  assign T318 = T319 - 1'h1;
  assign T319 = 1'h1 << T320;
  assign T320 = T321 + 2'h1;
  assign T321 = oacq_data_cnt - oacq_data_cnt;
  assign T322 = iacq_data_valid >> oacq_data_cnt;
  assign T422 = reset ? 4'h0 : T323;
  assign T323 = T59 ? T331 : T324;
  assign T324 = T229 ? T325 : iacq_data_valid;
  assign T325 = T329 | T326;
  assign T326 = T423 & T327;
  assign T327 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T423 = T328 ? 4'hf : 4'h0;
  assign T328 = 1'h1;
  assign T329 = iacq_data_valid & T330;
  assign T330 = ~ T327;
  assign T331 = T332 << io_inner_acquire_bits_addr_beat;
  assign T332 = io_inner_acquire_bits_is_builtin_type & T333;
  assign T333 = T335 | T334;
  assign T334 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T335 = T337 | T336;
  assign T336 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T337 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T338 = collect_iacq_data ^ 1'h1;
  assign T339 = pending_ognt_ack ^ 1'h1;
  assign T340 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T341;
  assign T341 = T102 ? T342 : 1'h0;
  assign T342 = T343 | io_outer_acquire_ready;
  assign T343 = T344 ^ 1'h1;
  assign T344 = T346 | T345;
  assign T345 = 3'h2 == io_inner_release_bits_r_type;
  assign T346 = T348 | T347;
  assign T347 = 3'h1 == io_inner_release_bits_r_type;
  assign T348 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T349;
  assign T349 = T424;
  assign T424 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T356;
  assign T356 = T357;
  assign T357 = xact_is_builtin_type ? T362 : T358;
  assign T358 = T361 ? 2'h1 : T359;
  assign T359 = T360 ? 2'h0 : 2'h2;
  assign T360 = xact_a_type == 3'h1;
  assign T361 = xact_a_type == 3'h0;
  assign T362 = T371 ? 2'h2 : T363;
  assign T363 = T370 ? 2'h0 : T364;
  assign T364 = T369 ? 2'h2 : T365;
  assign T365 = T368 ? 2'h0 : T366;
  assign T366 = T367 ? 2'h0 : 2'h2;
  assign T367 = xact_a_type == 3'h4;
  assign T368 = xact_a_type == 3'h2;
  assign T369 = xact_a_type == 3'h0;
  assign T370 = xact_a_type == 3'h3;
  assign T371 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T372;
  assign T372 = xact_addr_block;
  assign io_inner_probe_valid = T373;
  assign T373 = T102 ? T374 : 1'h0;
  assign T374 = pending_probes != 1'h0;
  assign T425 = T426[1'h0:1'h0];
  assign T426 = reset ? 4'h0 : T350;
  assign T350 = T355 ? T428 : T351;
  assign T351 = T91 ? mask_incoherent : T427;
  assign T427 = {3'h0, pending_probes};
  assign T428 = {2'h0, T352};
  assign T352 = T429 & T353;
  assign T353 = ~ T354;
  assign T354 = 1'h1 << 1'h0;
  assign T429 = {1'h0, pending_probes};
  assign T355 = T102 & io_inner_probe_ready;
  assign io_inner_finish_ready = T150;
  assign io_inner_grant_bits_client_id = T375;
  assign T375 = xact_client_id;
  assign io_inner_grant_bits_data = T376;
  assign T376 = 4'h0;
  assign io_inner_grant_bits_g_type = T377;
  assign T377 = T430;
  assign T430 = {1'h0, T378};
  assign T378 = xact_is_builtin_type ? T381 : T431;
  assign T431 = {1'h0, T379};
  assign T379 = T380 ? 2'h0 : 2'h1;
  assign T380 = xact_a_type == 3'h0;
  assign T381 = T392 ? 3'h4 : T382;
  assign T382 = T391 ? 3'h5 : T383;
  assign T383 = T390 ? 3'h3 : T384;
  assign T384 = T389 ? 3'h3 : T385;
  assign T385 = T388 ? 3'h4 : T386;
  assign T386 = T387 ? 3'h1 : 3'h3;
  assign T387 = xact_a_type == 3'h5;
  assign T388 = xact_a_type == 3'h4;
  assign T389 = xact_a_type == 3'h3;
  assign T390 = xact_a_type == 3'h2;
  assign T391 = xact_a_type == 3'h1;
  assign T392 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T393;
  assign T393 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T394;
  assign T394 = 4'h5;
  assign io_inner_grant_bits_client_xact_id = T395;
  assign T395 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T396;
  assign T396 = 2'h0;
  assign io_inner_grant_valid = T397;
  assign T397 = T148 ? 1'h1 : T398;
  assign T398 = T142 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T399;
  assign T399 = T60 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T185 <= 1'b1;
  if(!T186 && T185 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T175 <= 1'b1;
  if(!T176 && T175 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T151 <= 1'b1;
  if(!T152 && T151 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= 3'h0;
    end else if(T147) begin
      state <= T143;
    end else if(T129) begin
      state <= T125;
    end else if(T122) begin
      state <= 3'h5;
    end else if(T120) begin
      state <= T119;
    end else if(T117) begin
      state <= T115;
    end else if(T76) begin
      state <= T61;
    end else if(T59) begin
      state <= T19;
    end
    if(T59) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T59) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T406;
    if(reset) begin
      R107 <= 2'h0;
    end else if(T110) begin
      R107 <= T109;
    end
    if(reset) begin
      R133 <= 2'h0;
    end else if(T136) begin
      R133 <= T135;
    end
    if(T59) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T59) begin
      collect_iacq_data <= T172;
    end else if(T162) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R166 <= 2'h0;
    end else if(T169) begin
      R166 <= T168;
    end
    if(T59) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T59) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T120) begin
      pending_ognt_ack <= 1'h1;
    end else if(T103) begin
      pending_ognt_ack <= 1'h1;
    end else if(T211) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T230) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T225) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T238) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T236) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T247) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T245) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T253) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T251) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T59) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T59) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T59) begin
      iacq_data_valid <= T331;
    end else if(T229) begin
      iacq_data_valid <= T325;
    end
    pending_probes <= T425;
  end
endmodule

module BroadcastAcquireTracker_5(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T400;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T401;
  wire[2:0] T25;
  wire[2:0] T402;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire pending_outer_write_;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[3:0] mask_incoherent;
  wire[3:0] T403;
  wire T51;
  wire T52;
  wire[3:0] mask_self;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T404;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T405;
  wire T58;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[2:0] T62;
  wire pending_outer_read;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire pending_outer_write;
  wire T69;
  wire T70;
  reg [2:0] xact_a_type;
  wire[2:0] T71;
  wire T72;
  wire T73;
  wire T74;
  reg  xact_is_builtin_type;
  wire T75;
  wire T76;
  wire T77;
  reg  release_count;
  wire T406;
  wire[2:0] T407;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T408;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire T85;
  wire[1:0] T409;
  wire T86;
  wire[2:0] T410;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T411;
  wire T90;
  wire T91;
  wire[2:0] T412;
  wire T92;
  wire[2:0] T413;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire oacq_data_done;
  wire T104;
  wire T105;
  wire T106;
  reg [1:0] R107;
  wire[1:0] T414;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire[2:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire ignt_data_done;
  wire T130;
  wire T131;
  wire T132;
  reg [1:0] R133;
  wire[1:0] T415;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire[2:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  reg[0:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire T159;
  reg  collect_iacq_data;
  wire T416;
  wire T160;
  wire T161;
  wire T162;
  wire iacq_data_done;
  wire T163;
  wire T164;
  wire T165;
  reg [1:0] R166;
  wire[1:0] T417;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  reg[0:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  reg [1:0] xact_client_id;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  reg[0:0] T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  reg [25:0] xact_addr_block;
  wire[25:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  reg  pending_ognt_ack;
  wire T418;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[3:0] T214;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[3:0] T220;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T221;
  wire[3:0] T222;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T223;
  wire[3:0] T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[1:0] T228;
  wire T229;
  wire T230;
  wire T231;
  wire[3:0] T232;
  wire[1:0] T233;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T234;
  wire[3:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[1:0] T241;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T242;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T243;
  wire[3:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T249;
  wire[3:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] oacq_write_beat_data;
  wire T257;
  wire[3:0] oacq_probe_data;
  wire T258;
  wire[16:0] T259;
  wire[16:0] T260;
  wire[16:0] T261;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T419;
  wire[12:0] T262;
  wire[6:0] T263;
  wire[2:0] T264;
  reg [16:0] xact_union;
  wire[16:0] T265;
  wire[3:0] T266;
  wire[16:0] T267;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T268;
  wire[15:0] T269;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T270;
  wire[15:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[15:0] T279;
  wire[15:0] T280;
  wire[7:0] T281;
  wire[7:0] T420;
  wire T282;
  wire[1:0] T283;
  wire T284;
  wire[3:0] T285;
  wire[7:0] T286;
  wire[7:0] T421;
  wire T287;
  wire T288;
  wire T289;
  wire[16:0] oacq_probe_union;
  wire[16:0] T290;
  wire[15:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[2:0] T294;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T295;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T296;
  wire T297;
  wire T298;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T299;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T303;
  wire[1:0] T304;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T308;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T309;
  wire[25:0] T310;
  wire[25:0] T311;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T312;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire[1:0] T321;
  wire T322;
  reg [3:0] iacq_data_valid;
  wire[3:0] T422;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[3:0] T326;
  wire[3:0] T327;
  wire[3:0] T423;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire[1:0] T349;
  wire[1:0] T424;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[1:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[25:0] T372;
  wire T373;
  wire T374;
  reg  pending_probes;
  wire T425;
  wire[3:0] T426;
  wire[3:0] T350;
  wire[3:0] T351;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[1:0] T352;
  wire T353;
  wire T354;
  wire[1:0] T429;
  wire T355;
  wire[1:0] T375;
  wire[3:0] T376;
  wire[3:0] T377;
  wire[3:0] T430;
  wire[2:0] T378;
  wire[2:0] T431;
  wire[1:0] T379;
  wire T380;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] T384;
  wire[2:0] T385;
  wire[2:0] T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[3:0] T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire T397;
  wire T398;
  wire T399;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R107 = {1{$random}};
    R133 = {1{$random}};
    T151 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R166 = {1{$random}};
    T175 = 1'b0;
    xact_client_id = {1{$random}};
    T185 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T400 = reset ? 3'h0 : T11;
  assign T11 = T149 ? 3'h0 : T12;
  assign T12 = T147 ? T143 : T13;
  assign T13 = T129 ? T125 : T14;
  assign T14 = T122 ? 3'h5 : T15;
  assign T15 = T120 ? T119 : T16;
  assign T16 = T117 ? T115 : T17;
  assign T17 = T76 ? T61 : T18;
  assign T18 = T59 ? T19 : state;
  assign T19 = T50 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T44 ? T41 : T22;
  assign T22 = T40 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T401;
  assign T401 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T402;
  assign T402 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T39 ? 3'h4 : T29;
  assign T29 = T38 ? 3'h5 : T30;
  assign T30 = T37 ? 3'h3 : T31;
  assign T31 = T36 ? 3'h3 : T32;
  assign T32 = T35 ? 3'h4 : T33;
  assign T33 = T34 ? 3'h1 : 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h5;
  assign T35 = io_inner_acquire_bits_a_type == 3'h4;
  assign T36 = io_inner_acquire_bits_a_type == 3'h3;
  assign T37 = io_inner_acquire_bits_a_type == 3'h2;
  assign T38 = io_inner_acquire_bits_a_type == 3'h1;
  assign T39 = io_inner_acquire_bits_a_type == 3'h0;
  assign T40 = 4'h0 == T24;
  assign T41 = T43 | T42;
  assign T42 = 4'h4 == T24;
  assign T43 = 4'h5 == T24;
  assign T44 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T45;
  assign T45 = T47 | T46;
  assign T46 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T49 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T50 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T403;
  assign T403 = {3'h0, T51};
  assign T51 = ~ T52;
  assign T52 = io_incoherent_0;
  assign mask_self = T56 | T53;
  assign T53 = T404 & T54;
  assign T54 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T404 = T55 ? 4'hf : 4'h0;
  assign T55 = 1'h0;
  assign T56 = T405 & T57;
  assign T57 = ~ T54;
  assign T405 = {3'h0, T58};
  assign T58 = 1'h1;
  assign T59 = T60 & io_inner_acquire_valid;
  assign T60 = 3'h0 == state;
  assign T61 = pending_outer_write ? 3'h3 : T62;
  assign T62 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T66 : T63;
  assign T63 = T65 | T64;
  assign T64 = 4'h1 == io_inner_grant_bits_g_type;
  assign T65 = 4'h0 == io_inner_grant_bits_g_type;
  assign T66 = T68 | T67;
  assign T67 = 4'h4 == io_inner_grant_bits_g_type;
  assign T68 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T69;
  assign T69 = T72 | T70;
  assign T70 = 3'h4 == xact_a_type;
  assign T71 = T59 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T72 = T74 | T73;
  assign T73 = 3'h3 == xact_a_type;
  assign T74 = 3'h2 == xact_a_type;
  assign T75 = T59 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T76 = T103 & T77;
  assign T77 = release_count == 1'h1;
  assign T406 = T407[1'h0:1'h0];
  assign T407 = reset ? 3'h0 : T78;
  assign T78 = T94 ? T413 : T79;
  assign T79 = T103 ? T412 : T80;
  assign T80 = T91 ? T81 : T408;
  assign T408 = {2'h0, release_count};
  assign T81 = T410 + T82;
  assign T82 = {1'h0, T83};
  assign T83 = T409 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = mask_incoherent[2'h3:2'h3];
  assign T409 = {1'h0, T86};
  assign T86 = mask_incoherent[2'h2:2'h2];
  assign T410 = {1'h0, T87};
  assign T87 = T411 + T88;
  assign T88 = {1'h0, T89};
  assign T89 = mask_incoherent[1'h1:1'h1];
  assign T411 = {1'h0, T90};
  assign T90 = mask_incoherent[1'h0:1'h0];
  assign T91 = T59 & T50;
  assign T412 = {2'h0, T92};
  assign T92 = release_count - 1'h1;
  assign T413 = {2'h0, T93};
  assign T93 = release_count - 1'h1;
  assign T94 = T101 & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = T98 | T97;
  assign T97 = 3'h2 == io_inner_release_bits_r_type;
  assign T98 = T100 | T99;
  assign T99 = 3'h1 == io_inner_release_bits_r_type;
  assign T100 = 3'h0 == io_inner_release_bits_r_type;
  assign T101 = T102 & io_inner_release_valid;
  assign T102 = 3'h1 == state;
  assign T103 = T113 & oacq_data_done;
  assign oacq_data_done = T111 ? T105 : T104;
  assign T104 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T105 = T110 & T106;
  assign T106 = R107 == 2'h3;
  assign T414 = reset ? 2'h0 : T108;
  assign T108 = T110 ? T109 : R107;
  assign T109 = R107 + 2'h1;
  assign T110 = T104 & T111;
  assign T111 = io_outer_acquire_bits_is_builtin_type & T112;
  assign T112 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T113 = T114 & io_outer_acquire_ready;
  assign T114 = T101 & T96;
  assign T115 = pending_outer_write ? 3'h3 : T116;
  assign T116 = pending_outer_read ? 3'h2 : 3'h4;
  assign T117 = T94 & T118;
  assign T118 = release_count == 1'h1;
  assign T119 = pending_outer_read ? 3'h2 : 3'h5;
  assign T120 = T121 & oacq_data_done;
  assign T121 = 3'h3 == state;
  assign T122 = T124 & T123;
  assign T123 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T124 = 3'h2 == state;
  assign T125 = T126 ? 3'h6 : 3'h0;
  assign T126 = T127 ^ 1'h1;
  assign T127 = io_inner_grant_bits_is_builtin_type & T128;
  assign T128 = io_inner_grant_bits_g_type == 4'h0;
  assign T129 = T142 & ignt_data_done;
  assign ignt_data_done = T137 ? T131 : T130;
  assign T130 = io_inner_grant_ready & io_inner_grant_valid;
  assign T131 = T136 & T132;
  assign T132 = R133 == 2'h3;
  assign T415 = reset ? 2'h0 : T134;
  assign T134 = T136 ? T135 : R133;
  assign T135 = R133 + 2'h1;
  assign T136 = T130 & T137;
  assign T137 = io_inner_grant_bits_is_builtin_type ? T141 : T138;
  assign T138 = T140 | T139;
  assign T139 = 4'h1 == io_inner_grant_bits_g_type;
  assign T140 = 4'h0 == io_inner_grant_bits_g_type;
  assign T141 = 4'h5 == io_inner_grant_bits_g_type;
  assign T142 = 3'h5 == state;
  assign T143 = T144 ? 3'h6 : 3'h0;
  assign T144 = T145 ^ 1'h1;
  assign T145 = io_inner_grant_bits_is_builtin_type & T146;
  assign T146 = io_inner_grant_bits_g_type == 4'h0;
  assign T147 = T148 & io_inner_grant_ready;
  assign T148 = 3'h4 == state;
  assign T149 = T150 & io_inner_finish_valid;
  assign T150 = 3'h6 == state;
  assign T152 = T153 | reset;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T157 & T155;
  assign T155 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T156 = T59 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T157 = T159 & T158;
  assign T158 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T159 = T174 & collect_iacq_data;
  assign T416 = reset ? 1'h0 : T160;
  assign T160 = T59 ? T172 : T161;
  assign T161 = T162 ? 1'h0 : collect_iacq_data;
  assign T162 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T170 ? T164 : T163;
  assign T163 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T164 = T169 & T165;
  assign T165 = R166 == 2'h3;
  assign T417 = reset ? 2'h0 : T167;
  assign T167 = T169 ? T168 : R166;
  assign T168 = R166 + 2'h1;
  assign T169 = T163 & T170;
  assign T170 = io_inner_acquire_bits_is_builtin_type & T171;
  assign T171 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = state != 3'h0;
  assign T176 = T177 | reset;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T181 & T179;
  assign T179 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T180 = T59 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T181 = T183 & T182;
  assign T182 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T183 = T184 & collect_iacq_data;
  assign T184 = state != 3'h0;
  assign T186 = T187 | reset;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T192 & T189;
  assign T189 = T191 | T190;
  assign T190 = 3'h5 == xact_a_type;
  assign T191 = 3'h4 == xact_a_type;
  assign T192 = T193 & xact_is_builtin_type;
  assign T193 = state != 3'h0;
  assign io_has_release_match = T194;
  assign T194 = T196 & T195;
  assign T195 = state == 3'h1;
  assign T196 = T198 & T197;
  assign T197 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T198 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T199 = T59 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T200;
  assign T200 = T201 & collect_iacq_data;
  assign T201 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T202;
  assign T202 = T204 & T203;
  assign T203 = collect_iacq_data ^ 1'h1;
  assign T204 = T206 & T205;
  assign T205 = state != 3'h0;
  assign T206 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T207;
  assign T207 = T142 ? io_inner_grant_ready : pending_ognt_ack;
  assign T418 = reset ? 1'h0 : T208;
  assign T208 = T120 ? 1'h1 : T209;
  assign T209 = T103 ? 1'h1 : T210;
  assign T210 = T211 ? 1'h0 : pending_ognt_ack;
  assign T211 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T212;
  assign T212 = T258 ? oacq_probe_data : T213;
  assign T213 = T257 ? T220 : T214;
  assign T214 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T215;
  assign T215 = T217 | T216;
  assign T216 = 3'h4 == xact_a_type;
  assign T217 = T219 | T218;
  assign T218 = 3'h0 == xact_a_type;
  assign T219 = 3'h2 == xact_a_type;
  assign T220 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T221;
  assign T221 = T256 ? T242 : T222;
  assign T222 = T240 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T223 = T230 ? io_inner_acquire_bits_data : T224;
  assign T224 = T225 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T225 = T229 & T226;
  assign T226 = T227[1'h0:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = io_inner_acquire_bits_addr_beat;
  assign T229 = collect_iacq_data & io_inner_acquire_valid;
  assign T230 = T59 & T231;
  assign T231 = T232[1'h0:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = 2'h0;
  assign T234 = T238 ? io_inner_acquire_bits_data : T235;
  assign T235 = T236 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T236 = T229 & T237;
  assign T237 = T227[1'h1:1'h1];
  assign T238 = T59 & T239;
  assign T239 = T232[1'h1:1'h1];
  assign T240 = T241[1'h0:1'h0];
  assign T241 = oacq_data_cnt;
  assign oacq_data_cnt = T111 ? R107 : 2'h0;
  assign T242 = T255 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T243 = T247 ? io_inner_acquire_bits_data : T244;
  assign T244 = T245 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T245 = T229 & T246;
  assign T246 = T227[2'h2:2'h2];
  assign T247 = T59 & T248;
  assign T248 = T232[2'h2:2'h2];
  assign T249 = T253 ? io_inner_acquire_bits_data : T250;
  assign T250 = T251 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T251 = T229 & T252;
  assign T252 = T227[2'h3:2'h3];
  assign T253 = T59 & T254;
  assign T254 = T232[2'h3:2'h3];
  assign T255 = T241[1'h0:1'h0];
  assign T256 = T241[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T257 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T258 = state == 3'h1;
  assign io_outer_acquire_bits_union = T259;
  assign T259 = T258 ? oacq_probe_union : T260;
  assign T260 = T257 ? T267 : T261;
  assign T261 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T419;
  assign T419 = {4'h0, T262};
  assign T262 = {T263, 6'h0};
  assign T263 = {T266, T264};
  assign T264 = xact_union[4'h8:3'h6];
  assign T265 = T59 ? io_inner_acquire_bits_union : xact_union;
  assign T266 = xact_union[4'hc:4'h9];
  assign T267 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T268;
  assign T268 = {T269, 1'h1};
  assign T269 = 16'hffff;
  assign oacq_write_beat_union = T270;
  assign T270 = {T271, 1'h1};
  assign T271 = T288 ? T279 : T272;
  assign T272 = T274 ? T273 : 16'h0;
  assign T273 = xact_union[5'h10:1'h1];
  assign T274 = T277 | T275;
  assign T275 = xact_is_builtin_type & T276;
  assign T276 = xact_a_type == 3'h2;
  assign T277 = xact_is_builtin_type & T278;
  assign T278 = xact_a_type == 3'h3;
  assign T279 = T280;
  assign T280 = {T286, T281};
  assign T281 = 8'h0 - T420;
  assign T420 = {7'h0, T282};
  assign T282 = T283[1'h0:1'h0];
  assign T283 = 1'h1 << T284;
  assign T284 = T285[2'h3:2'h3];
  assign T285 = xact_union[4'hc:4'h9];
  assign T286 = 8'h0 - T421;
  assign T421 = {7'h0, T287};
  assign T287 = T283[1'h1:1'h1];
  assign T288 = xact_is_builtin_type & T289;
  assign T289 = xact_a_type == 3'h4;
  assign oacq_probe_union = T290;
  assign T290 = {T291, 1'h1};
  assign T291 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T292;
  assign T292 = T258 ? oacq_probe_a_type : T293;
  assign T293 = T257 ? T295 : T294;
  assign T294 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T295 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T296;
  assign T296 = T258 ? oacq_probe_is_builtin_type : T297;
  assign T297 = T257 ? T299 : T298;
  assign T298 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T299 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T300;
  assign T300 = T258 ? oacq_probe_addr_beat : T301;
  assign T301 = T257 ? T304 : T302;
  assign T302 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T303 = T59 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T304 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T305;
  assign T305 = T258 ? oacq_probe_client_xact_id : T306;
  assign T306 = T257 ? T308 : T307;
  assign T307 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h6;
  assign oacq_read_beat_client_xact_id = 4'h6;
  assign T308 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h6;
  assign oacq_write_beat_client_xact_id = 4'h6;
  assign oacq_probe_client_xact_id = 4'h6;
  assign io_outer_acquire_bits_addr_block = T309;
  assign T309 = T258 ? oacq_probe_addr_block : T310;
  assign T310 = T257 ? T312 : T311;
  assign T311 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T312 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T313;
  assign T313 = T124 ? T340 : T314;
  assign T314 = T121 ? T315 : T114;
  assign T315 = T339 & T316;
  assign T316 = T338 | T317;
  assign T317 = T322 & T318;
  assign T318 = T319 - 1'h1;
  assign T319 = 1'h1 << T320;
  assign T320 = T321 + 2'h1;
  assign T321 = oacq_data_cnt - oacq_data_cnt;
  assign T322 = iacq_data_valid >> oacq_data_cnt;
  assign T422 = reset ? 4'h0 : T323;
  assign T323 = T59 ? T331 : T324;
  assign T324 = T229 ? T325 : iacq_data_valid;
  assign T325 = T329 | T326;
  assign T326 = T423 & T327;
  assign T327 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T423 = T328 ? 4'hf : 4'h0;
  assign T328 = 1'h1;
  assign T329 = iacq_data_valid & T330;
  assign T330 = ~ T327;
  assign T331 = T332 << io_inner_acquire_bits_addr_beat;
  assign T332 = io_inner_acquire_bits_is_builtin_type & T333;
  assign T333 = T335 | T334;
  assign T334 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T335 = T337 | T336;
  assign T336 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T337 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T338 = collect_iacq_data ^ 1'h1;
  assign T339 = pending_ognt_ack ^ 1'h1;
  assign T340 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T341;
  assign T341 = T102 ? T342 : 1'h0;
  assign T342 = T343 | io_outer_acquire_ready;
  assign T343 = T344 ^ 1'h1;
  assign T344 = T346 | T345;
  assign T345 = 3'h2 == io_inner_release_bits_r_type;
  assign T346 = T348 | T347;
  assign T347 = 3'h1 == io_inner_release_bits_r_type;
  assign T348 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T349;
  assign T349 = T424;
  assign T424 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T356;
  assign T356 = T357;
  assign T357 = xact_is_builtin_type ? T362 : T358;
  assign T358 = T361 ? 2'h1 : T359;
  assign T359 = T360 ? 2'h0 : 2'h2;
  assign T360 = xact_a_type == 3'h1;
  assign T361 = xact_a_type == 3'h0;
  assign T362 = T371 ? 2'h2 : T363;
  assign T363 = T370 ? 2'h0 : T364;
  assign T364 = T369 ? 2'h2 : T365;
  assign T365 = T368 ? 2'h0 : T366;
  assign T366 = T367 ? 2'h0 : 2'h2;
  assign T367 = xact_a_type == 3'h4;
  assign T368 = xact_a_type == 3'h2;
  assign T369 = xact_a_type == 3'h0;
  assign T370 = xact_a_type == 3'h3;
  assign T371 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T372;
  assign T372 = xact_addr_block;
  assign io_inner_probe_valid = T373;
  assign T373 = T102 ? T374 : 1'h0;
  assign T374 = pending_probes != 1'h0;
  assign T425 = T426[1'h0:1'h0];
  assign T426 = reset ? 4'h0 : T350;
  assign T350 = T355 ? T428 : T351;
  assign T351 = T91 ? mask_incoherent : T427;
  assign T427 = {3'h0, pending_probes};
  assign T428 = {2'h0, T352};
  assign T352 = T429 & T353;
  assign T353 = ~ T354;
  assign T354 = 1'h1 << 1'h0;
  assign T429 = {1'h0, pending_probes};
  assign T355 = T102 & io_inner_probe_ready;
  assign io_inner_finish_ready = T150;
  assign io_inner_grant_bits_client_id = T375;
  assign T375 = xact_client_id;
  assign io_inner_grant_bits_data = T376;
  assign T376 = 4'h0;
  assign io_inner_grant_bits_g_type = T377;
  assign T377 = T430;
  assign T430 = {1'h0, T378};
  assign T378 = xact_is_builtin_type ? T381 : T431;
  assign T431 = {1'h0, T379};
  assign T379 = T380 ? 2'h0 : 2'h1;
  assign T380 = xact_a_type == 3'h0;
  assign T381 = T392 ? 3'h4 : T382;
  assign T382 = T391 ? 3'h5 : T383;
  assign T383 = T390 ? 3'h3 : T384;
  assign T384 = T389 ? 3'h3 : T385;
  assign T385 = T388 ? 3'h4 : T386;
  assign T386 = T387 ? 3'h1 : 3'h3;
  assign T387 = xact_a_type == 3'h5;
  assign T388 = xact_a_type == 3'h4;
  assign T389 = xact_a_type == 3'h3;
  assign T390 = xact_a_type == 3'h2;
  assign T391 = xact_a_type == 3'h1;
  assign T392 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T393;
  assign T393 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T394;
  assign T394 = 4'h6;
  assign io_inner_grant_bits_client_xact_id = T395;
  assign T395 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T396;
  assign T396 = 2'h0;
  assign io_inner_grant_valid = T397;
  assign T397 = T148 ? 1'h1 : T398;
  assign T398 = T142 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T399;
  assign T399 = T60 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T185 <= 1'b1;
  if(!T186 && T185 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T175 <= 1'b1;
  if(!T176 && T175 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T151 <= 1'b1;
  if(!T152 && T151 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= 3'h0;
    end else if(T147) begin
      state <= T143;
    end else if(T129) begin
      state <= T125;
    end else if(T122) begin
      state <= 3'h5;
    end else if(T120) begin
      state <= T119;
    end else if(T117) begin
      state <= T115;
    end else if(T76) begin
      state <= T61;
    end else if(T59) begin
      state <= T19;
    end
    if(T59) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T59) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T406;
    if(reset) begin
      R107 <= 2'h0;
    end else if(T110) begin
      R107 <= T109;
    end
    if(reset) begin
      R133 <= 2'h0;
    end else if(T136) begin
      R133 <= T135;
    end
    if(T59) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T59) begin
      collect_iacq_data <= T172;
    end else if(T162) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R166 <= 2'h0;
    end else if(T169) begin
      R166 <= T168;
    end
    if(T59) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T59) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T120) begin
      pending_ognt_ack <= 1'h1;
    end else if(T103) begin
      pending_ognt_ack <= 1'h1;
    end else if(T211) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T230) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T225) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T238) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T236) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T247) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T245) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T253) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T251) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T59) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T59) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T59) begin
      iacq_data_valid <= T331;
    end else if(T229) begin
      iacq_data_valid <= T325;
    end
    pending_probes <= T425;
  end
endmodule

module BroadcastAcquireTracker_6(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T400;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T401;
  wire[2:0] T25;
  wire[2:0] T402;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire pending_outer_write_;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[3:0] mask_incoherent;
  wire[3:0] T403;
  wire T51;
  wire T52;
  wire[3:0] mask_self;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T404;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T405;
  wire T58;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[2:0] T62;
  wire pending_outer_read;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire pending_outer_write;
  wire T69;
  wire T70;
  reg [2:0] xact_a_type;
  wire[2:0] T71;
  wire T72;
  wire T73;
  wire T74;
  reg  xact_is_builtin_type;
  wire T75;
  wire T76;
  wire T77;
  reg  release_count;
  wire T406;
  wire[2:0] T407;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T408;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire T85;
  wire[1:0] T409;
  wire T86;
  wire[2:0] T410;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T411;
  wire T90;
  wire T91;
  wire[2:0] T412;
  wire T92;
  wire[2:0] T413;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire oacq_data_done;
  wire T104;
  wire T105;
  wire T106;
  reg [1:0] R107;
  wire[1:0] T414;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire[2:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire ignt_data_done;
  wire T130;
  wire T131;
  wire T132;
  reg [1:0] R133;
  wire[1:0] T415;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire[2:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  reg[0:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire T159;
  reg  collect_iacq_data;
  wire T416;
  wire T160;
  wire T161;
  wire T162;
  wire iacq_data_done;
  wire T163;
  wire T164;
  wire T165;
  reg [1:0] R166;
  wire[1:0] T417;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  reg[0:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  reg [1:0] xact_client_id;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  reg[0:0] T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  reg [25:0] xact_addr_block;
  wire[25:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  reg  pending_ognt_ack;
  wire T418;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[3:0] T214;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[3:0] T220;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T221;
  wire[3:0] T222;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T223;
  wire[3:0] T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[1:0] T228;
  wire T229;
  wire T230;
  wire T231;
  wire[3:0] T232;
  wire[1:0] T233;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T234;
  wire[3:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[1:0] T241;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T242;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T243;
  wire[3:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T249;
  wire[3:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] oacq_write_beat_data;
  wire T257;
  wire[3:0] oacq_probe_data;
  wire T258;
  wire[16:0] T259;
  wire[16:0] T260;
  wire[16:0] T261;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T419;
  wire[12:0] T262;
  wire[6:0] T263;
  wire[2:0] T264;
  reg [16:0] xact_union;
  wire[16:0] T265;
  wire[3:0] T266;
  wire[16:0] T267;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T268;
  wire[15:0] T269;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T270;
  wire[15:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[15:0] T279;
  wire[15:0] T280;
  wire[7:0] T281;
  wire[7:0] T420;
  wire T282;
  wire[1:0] T283;
  wire T284;
  wire[3:0] T285;
  wire[7:0] T286;
  wire[7:0] T421;
  wire T287;
  wire T288;
  wire T289;
  wire[16:0] oacq_probe_union;
  wire[16:0] T290;
  wire[15:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[2:0] T294;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T295;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T296;
  wire T297;
  wire T298;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T299;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T303;
  wire[1:0] T304;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T308;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T309;
  wire[25:0] T310;
  wire[25:0] T311;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T312;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire[1:0] T321;
  wire T322;
  reg [3:0] iacq_data_valid;
  wire[3:0] T422;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[3:0] T326;
  wire[3:0] T327;
  wire[3:0] T423;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire[1:0] T349;
  wire[1:0] T424;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[1:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[25:0] T372;
  wire T373;
  wire T374;
  reg  pending_probes;
  wire T425;
  wire[3:0] T426;
  wire[3:0] T350;
  wire[3:0] T351;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[1:0] T352;
  wire T353;
  wire T354;
  wire[1:0] T429;
  wire T355;
  wire[1:0] T375;
  wire[3:0] T376;
  wire[3:0] T377;
  wire[3:0] T430;
  wire[2:0] T378;
  wire[2:0] T431;
  wire[1:0] T379;
  wire T380;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] T384;
  wire[2:0] T385;
  wire[2:0] T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[3:0] T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire T397;
  wire T398;
  wire T399;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R107 = {1{$random}};
    R133 = {1{$random}};
    T151 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R166 = {1{$random}};
    T175 = 1'b0;
    xact_client_id = {1{$random}};
    T185 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T400 = reset ? 3'h0 : T11;
  assign T11 = T149 ? 3'h0 : T12;
  assign T12 = T147 ? T143 : T13;
  assign T13 = T129 ? T125 : T14;
  assign T14 = T122 ? 3'h5 : T15;
  assign T15 = T120 ? T119 : T16;
  assign T16 = T117 ? T115 : T17;
  assign T17 = T76 ? T61 : T18;
  assign T18 = T59 ? T19 : state;
  assign T19 = T50 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T44 ? T41 : T22;
  assign T22 = T40 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T401;
  assign T401 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T402;
  assign T402 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T39 ? 3'h4 : T29;
  assign T29 = T38 ? 3'h5 : T30;
  assign T30 = T37 ? 3'h3 : T31;
  assign T31 = T36 ? 3'h3 : T32;
  assign T32 = T35 ? 3'h4 : T33;
  assign T33 = T34 ? 3'h1 : 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h5;
  assign T35 = io_inner_acquire_bits_a_type == 3'h4;
  assign T36 = io_inner_acquire_bits_a_type == 3'h3;
  assign T37 = io_inner_acquire_bits_a_type == 3'h2;
  assign T38 = io_inner_acquire_bits_a_type == 3'h1;
  assign T39 = io_inner_acquire_bits_a_type == 3'h0;
  assign T40 = 4'h0 == T24;
  assign T41 = T43 | T42;
  assign T42 = 4'h4 == T24;
  assign T43 = 4'h5 == T24;
  assign T44 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T45;
  assign T45 = T47 | T46;
  assign T46 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T49 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T50 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T403;
  assign T403 = {3'h0, T51};
  assign T51 = ~ T52;
  assign T52 = io_incoherent_0;
  assign mask_self = T56 | T53;
  assign T53 = T404 & T54;
  assign T54 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T404 = T55 ? 4'hf : 4'h0;
  assign T55 = 1'h0;
  assign T56 = T405 & T57;
  assign T57 = ~ T54;
  assign T405 = {3'h0, T58};
  assign T58 = 1'h1;
  assign T59 = T60 & io_inner_acquire_valid;
  assign T60 = 3'h0 == state;
  assign T61 = pending_outer_write ? 3'h3 : T62;
  assign T62 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T66 : T63;
  assign T63 = T65 | T64;
  assign T64 = 4'h1 == io_inner_grant_bits_g_type;
  assign T65 = 4'h0 == io_inner_grant_bits_g_type;
  assign T66 = T68 | T67;
  assign T67 = 4'h4 == io_inner_grant_bits_g_type;
  assign T68 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T69;
  assign T69 = T72 | T70;
  assign T70 = 3'h4 == xact_a_type;
  assign T71 = T59 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T72 = T74 | T73;
  assign T73 = 3'h3 == xact_a_type;
  assign T74 = 3'h2 == xact_a_type;
  assign T75 = T59 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T76 = T103 & T77;
  assign T77 = release_count == 1'h1;
  assign T406 = T407[1'h0:1'h0];
  assign T407 = reset ? 3'h0 : T78;
  assign T78 = T94 ? T413 : T79;
  assign T79 = T103 ? T412 : T80;
  assign T80 = T91 ? T81 : T408;
  assign T408 = {2'h0, release_count};
  assign T81 = T410 + T82;
  assign T82 = {1'h0, T83};
  assign T83 = T409 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = mask_incoherent[2'h3:2'h3];
  assign T409 = {1'h0, T86};
  assign T86 = mask_incoherent[2'h2:2'h2];
  assign T410 = {1'h0, T87};
  assign T87 = T411 + T88;
  assign T88 = {1'h0, T89};
  assign T89 = mask_incoherent[1'h1:1'h1];
  assign T411 = {1'h0, T90};
  assign T90 = mask_incoherent[1'h0:1'h0];
  assign T91 = T59 & T50;
  assign T412 = {2'h0, T92};
  assign T92 = release_count - 1'h1;
  assign T413 = {2'h0, T93};
  assign T93 = release_count - 1'h1;
  assign T94 = T101 & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = T98 | T97;
  assign T97 = 3'h2 == io_inner_release_bits_r_type;
  assign T98 = T100 | T99;
  assign T99 = 3'h1 == io_inner_release_bits_r_type;
  assign T100 = 3'h0 == io_inner_release_bits_r_type;
  assign T101 = T102 & io_inner_release_valid;
  assign T102 = 3'h1 == state;
  assign T103 = T113 & oacq_data_done;
  assign oacq_data_done = T111 ? T105 : T104;
  assign T104 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T105 = T110 & T106;
  assign T106 = R107 == 2'h3;
  assign T414 = reset ? 2'h0 : T108;
  assign T108 = T110 ? T109 : R107;
  assign T109 = R107 + 2'h1;
  assign T110 = T104 & T111;
  assign T111 = io_outer_acquire_bits_is_builtin_type & T112;
  assign T112 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T113 = T114 & io_outer_acquire_ready;
  assign T114 = T101 & T96;
  assign T115 = pending_outer_write ? 3'h3 : T116;
  assign T116 = pending_outer_read ? 3'h2 : 3'h4;
  assign T117 = T94 & T118;
  assign T118 = release_count == 1'h1;
  assign T119 = pending_outer_read ? 3'h2 : 3'h5;
  assign T120 = T121 & oacq_data_done;
  assign T121 = 3'h3 == state;
  assign T122 = T124 & T123;
  assign T123 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T124 = 3'h2 == state;
  assign T125 = T126 ? 3'h6 : 3'h0;
  assign T126 = T127 ^ 1'h1;
  assign T127 = io_inner_grant_bits_is_builtin_type & T128;
  assign T128 = io_inner_grant_bits_g_type == 4'h0;
  assign T129 = T142 & ignt_data_done;
  assign ignt_data_done = T137 ? T131 : T130;
  assign T130 = io_inner_grant_ready & io_inner_grant_valid;
  assign T131 = T136 & T132;
  assign T132 = R133 == 2'h3;
  assign T415 = reset ? 2'h0 : T134;
  assign T134 = T136 ? T135 : R133;
  assign T135 = R133 + 2'h1;
  assign T136 = T130 & T137;
  assign T137 = io_inner_grant_bits_is_builtin_type ? T141 : T138;
  assign T138 = T140 | T139;
  assign T139 = 4'h1 == io_inner_grant_bits_g_type;
  assign T140 = 4'h0 == io_inner_grant_bits_g_type;
  assign T141 = 4'h5 == io_inner_grant_bits_g_type;
  assign T142 = 3'h5 == state;
  assign T143 = T144 ? 3'h6 : 3'h0;
  assign T144 = T145 ^ 1'h1;
  assign T145 = io_inner_grant_bits_is_builtin_type & T146;
  assign T146 = io_inner_grant_bits_g_type == 4'h0;
  assign T147 = T148 & io_inner_grant_ready;
  assign T148 = 3'h4 == state;
  assign T149 = T150 & io_inner_finish_valid;
  assign T150 = 3'h6 == state;
  assign T152 = T153 | reset;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T157 & T155;
  assign T155 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T156 = T59 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T157 = T159 & T158;
  assign T158 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T159 = T174 & collect_iacq_data;
  assign T416 = reset ? 1'h0 : T160;
  assign T160 = T59 ? T172 : T161;
  assign T161 = T162 ? 1'h0 : collect_iacq_data;
  assign T162 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T170 ? T164 : T163;
  assign T163 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T164 = T169 & T165;
  assign T165 = R166 == 2'h3;
  assign T417 = reset ? 2'h0 : T167;
  assign T167 = T169 ? T168 : R166;
  assign T168 = R166 + 2'h1;
  assign T169 = T163 & T170;
  assign T170 = io_inner_acquire_bits_is_builtin_type & T171;
  assign T171 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = state != 3'h0;
  assign T176 = T177 | reset;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T181 & T179;
  assign T179 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T180 = T59 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T181 = T183 & T182;
  assign T182 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T183 = T184 & collect_iacq_data;
  assign T184 = state != 3'h0;
  assign T186 = T187 | reset;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T192 & T189;
  assign T189 = T191 | T190;
  assign T190 = 3'h5 == xact_a_type;
  assign T191 = 3'h4 == xact_a_type;
  assign T192 = T193 & xact_is_builtin_type;
  assign T193 = state != 3'h0;
  assign io_has_release_match = T194;
  assign T194 = T196 & T195;
  assign T195 = state == 3'h1;
  assign T196 = T198 & T197;
  assign T197 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T198 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T199 = T59 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T200;
  assign T200 = T201 & collect_iacq_data;
  assign T201 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T202;
  assign T202 = T204 & T203;
  assign T203 = collect_iacq_data ^ 1'h1;
  assign T204 = T206 & T205;
  assign T205 = state != 3'h0;
  assign T206 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T207;
  assign T207 = T142 ? io_inner_grant_ready : pending_ognt_ack;
  assign T418 = reset ? 1'h0 : T208;
  assign T208 = T120 ? 1'h1 : T209;
  assign T209 = T103 ? 1'h1 : T210;
  assign T210 = T211 ? 1'h0 : pending_ognt_ack;
  assign T211 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T212;
  assign T212 = T258 ? oacq_probe_data : T213;
  assign T213 = T257 ? T220 : T214;
  assign T214 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T215;
  assign T215 = T217 | T216;
  assign T216 = 3'h4 == xact_a_type;
  assign T217 = T219 | T218;
  assign T218 = 3'h0 == xact_a_type;
  assign T219 = 3'h2 == xact_a_type;
  assign T220 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T221;
  assign T221 = T256 ? T242 : T222;
  assign T222 = T240 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T223 = T230 ? io_inner_acquire_bits_data : T224;
  assign T224 = T225 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T225 = T229 & T226;
  assign T226 = T227[1'h0:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = io_inner_acquire_bits_addr_beat;
  assign T229 = collect_iacq_data & io_inner_acquire_valid;
  assign T230 = T59 & T231;
  assign T231 = T232[1'h0:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = 2'h0;
  assign T234 = T238 ? io_inner_acquire_bits_data : T235;
  assign T235 = T236 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T236 = T229 & T237;
  assign T237 = T227[1'h1:1'h1];
  assign T238 = T59 & T239;
  assign T239 = T232[1'h1:1'h1];
  assign T240 = T241[1'h0:1'h0];
  assign T241 = oacq_data_cnt;
  assign oacq_data_cnt = T111 ? R107 : 2'h0;
  assign T242 = T255 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T243 = T247 ? io_inner_acquire_bits_data : T244;
  assign T244 = T245 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T245 = T229 & T246;
  assign T246 = T227[2'h2:2'h2];
  assign T247 = T59 & T248;
  assign T248 = T232[2'h2:2'h2];
  assign T249 = T253 ? io_inner_acquire_bits_data : T250;
  assign T250 = T251 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T251 = T229 & T252;
  assign T252 = T227[2'h3:2'h3];
  assign T253 = T59 & T254;
  assign T254 = T232[2'h3:2'h3];
  assign T255 = T241[1'h0:1'h0];
  assign T256 = T241[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T257 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T258 = state == 3'h1;
  assign io_outer_acquire_bits_union = T259;
  assign T259 = T258 ? oacq_probe_union : T260;
  assign T260 = T257 ? T267 : T261;
  assign T261 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T419;
  assign T419 = {4'h0, T262};
  assign T262 = {T263, 6'h0};
  assign T263 = {T266, T264};
  assign T264 = xact_union[4'h8:3'h6];
  assign T265 = T59 ? io_inner_acquire_bits_union : xact_union;
  assign T266 = xact_union[4'hc:4'h9];
  assign T267 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T268;
  assign T268 = {T269, 1'h1};
  assign T269 = 16'hffff;
  assign oacq_write_beat_union = T270;
  assign T270 = {T271, 1'h1};
  assign T271 = T288 ? T279 : T272;
  assign T272 = T274 ? T273 : 16'h0;
  assign T273 = xact_union[5'h10:1'h1];
  assign T274 = T277 | T275;
  assign T275 = xact_is_builtin_type & T276;
  assign T276 = xact_a_type == 3'h2;
  assign T277 = xact_is_builtin_type & T278;
  assign T278 = xact_a_type == 3'h3;
  assign T279 = T280;
  assign T280 = {T286, T281};
  assign T281 = 8'h0 - T420;
  assign T420 = {7'h0, T282};
  assign T282 = T283[1'h0:1'h0];
  assign T283 = 1'h1 << T284;
  assign T284 = T285[2'h3:2'h3];
  assign T285 = xact_union[4'hc:4'h9];
  assign T286 = 8'h0 - T421;
  assign T421 = {7'h0, T287};
  assign T287 = T283[1'h1:1'h1];
  assign T288 = xact_is_builtin_type & T289;
  assign T289 = xact_a_type == 3'h4;
  assign oacq_probe_union = T290;
  assign T290 = {T291, 1'h1};
  assign T291 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T292;
  assign T292 = T258 ? oacq_probe_a_type : T293;
  assign T293 = T257 ? T295 : T294;
  assign T294 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T295 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T296;
  assign T296 = T258 ? oacq_probe_is_builtin_type : T297;
  assign T297 = T257 ? T299 : T298;
  assign T298 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T299 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T300;
  assign T300 = T258 ? oacq_probe_addr_beat : T301;
  assign T301 = T257 ? T304 : T302;
  assign T302 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T303 = T59 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T304 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T305;
  assign T305 = T258 ? oacq_probe_client_xact_id : T306;
  assign T306 = T257 ? T308 : T307;
  assign T307 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h7;
  assign oacq_read_beat_client_xact_id = 4'h7;
  assign T308 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h7;
  assign oacq_write_beat_client_xact_id = 4'h7;
  assign oacq_probe_client_xact_id = 4'h7;
  assign io_outer_acquire_bits_addr_block = T309;
  assign T309 = T258 ? oacq_probe_addr_block : T310;
  assign T310 = T257 ? T312 : T311;
  assign T311 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T312 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T313;
  assign T313 = T124 ? T340 : T314;
  assign T314 = T121 ? T315 : T114;
  assign T315 = T339 & T316;
  assign T316 = T338 | T317;
  assign T317 = T322 & T318;
  assign T318 = T319 - 1'h1;
  assign T319 = 1'h1 << T320;
  assign T320 = T321 + 2'h1;
  assign T321 = oacq_data_cnt - oacq_data_cnt;
  assign T322 = iacq_data_valid >> oacq_data_cnt;
  assign T422 = reset ? 4'h0 : T323;
  assign T323 = T59 ? T331 : T324;
  assign T324 = T229 ? T325 : iacq_data_valid;
  assign T325 = T329 | T326;
  assign T326 = T423 & T327;
  assign T327 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T423 = T328 ? 4'hf : 4'h0;
  assign T328 = 1'h1;
  assign T329 = iacq_data_valid & T330;
  assign T330 = ~ T327;
  assign T331 = T332 << io_inner_acquire_bits_addr_beat;
  assign T332 = io_inner_acquire_bits_is_builtin_type & T333;
  assign T333 = T335 | T334;
  assign T334 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T335 = T337 | T336;
  assign T336 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T337 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T338 = collect_iacq_data ^ 1'h1;
  assign T339 = pending_ognt_ack ^ 1'h1;
  assign T340 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T341;
  assign T341 = T102 ? T342 : 1'h0;
  assign T342 = T343 | io_outer_acquire_ready;
  assign T343 = T344 ^ 1'h1;
  assign T344 = T346 | T345;
  assign T345 = 3'h2 == io_inner_release_bits_r_type;
  assign T346 = T348 | T347;
  assign T347 = 3'h1 == io_inner_release_bits_r_type;
  assign T348 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T349;
  assign T349 = T424;
  assign T424 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T356;
  assign T356 = T357;
  assign T357 = xact_is_builtin_type ? T362 : T358;
  assign T358 = T361 ? 2'h1 : T359;
  assign T359 = T360 ? 2'h0 : 2'h2;
  assign T360 = xact_a_type == 3'h1;
  assign T361 = xact_a_type == 3'h0;
  assign T362 = T371 ? 2'h2 : T363;
  assign T363 = T370 ? 2'h0 : T364;
  assign T364 = T369 ? 2'h2 : T365;
  assign T365 = T368 ? 2'h0 : T366;
  assign T366 = T367 ? 2'h0 : 2'h2;
  assign T367 = xact_a_type == 3'h4;
  assign T368 = xact_a_type == 3'h2;
  assign T369 = xact_a_type == 3'h0;
  assign T370 = xact_a_type == 3'h3;
  assign T371 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T372;
  assign T372 = xact_addr_block;
  assign io_inner_probe_valid = T373;
  assign T373 = T102 ? T374 : 1'h0;
  assign T374 = pending_probes != 1'h0;
  assign T425 = T426[1'h0:1'h0];
  assign T426 = reset ? 4'h0 : T350;
  assign T350 = T355 ? T428 : T351;
  assign T351 = T91 ? mask_incoherent : T427;
  assign T427 = {3'h0, pending_probes};
  assign T428 = {2'h0, T352};
  assign T352 = T429 & T353;
  assign T353 = ~ T354;
  assign T354 = 1'h1 << 1'h0;
  assign T429 = {1'h0, pending_probes};
  assign T355 = T102 & io_inner_probe_ready;
  assign io_inner_finish_ready = T150;
  assign io_inner_grant_bits_client_id = T375;
  assign T375 = xact_client_id;
  assign io_inner_grant_bits_data = T376;
  assign T376 = 4'h0;
  assign io_inner_grant_bits_g_type = T377;
  assign T377 = T430;
  assign T430 = {1'h0, T378};
  assign T378 = xact_is_builtin_type ? T381 : T431;
  assign T431 = {1'h0, T379};
  assign T379 = T380 ? 2'h0 : 2'h1;
  assign T380 = xact_a_type == 3'h0;
  assign T381 = T392 ? 3'h4 : T382;
  assign T382 = T391 ? 3'h5 : T383;
  assign T383 = T390 ? 3'h3 : T384;
  assign T384 = T389 ? 3'h3 : T385;
  assign T385 = T388 ? 3'h4 : T386;
  assign T386 = T387 ? 3'h1 : 3'h3;
  assign T387 = xact_a_type == 3'h5;
  assign T388 = xact_a_type == 3'h4;
  assign T389 = xact_a_type == 3'h3;
  assign T390 = xact_a_type == 3'h2;
  assign T391 = xact_a_type == 3'h1;
  assign T392 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T393;
  assign T393 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T394;
  assign T394 = 4'h7;
  assign io_inner_grant_bits_client_xact_id = T395;
  assign T395 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T396;
  assign T396 = 2'h0;
  assign io_inner_grant_valid = T397;
  assign T397 = T148 ? 1'h1 : T398;
  assign T398 = T142 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T399;
  assign T399 = T60 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T185 <= 1'b1;
  if(!T186 && T185 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T175 <= 1'b1;
  if(!T176 && T175 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T151 <= 1'b1;
  if(!T152 && T151 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= 3'h0;
    end else if(T147) begin
      state <= T143;
    end else if(T129) begin
      state <= T125;
    end else if(T122) begin
      state <= 3'h5;
    end else if(T120) begin
      state <= T119;
    end else if(T117) begin
      state <= T115;
    end else if(T76) begin
      state <= T61;
    end else if(T59) begin
      state <= T19;
    end
    if(T59) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T59) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T406;
    if(reset) begin
      R107 <= 2'h0;
    end else if(T110) begin
      R107 <= T109;
    end
    if(reset) begin
      R133 <= 2'h0;
    end else if(T136) begin
      R133 <= T135;
    end
    if(T59) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T59) begin
      collect_iacq_data <= T172;
    end else if(T162) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R166 <= 2'h0;
    end else if(T169) begin
      R166 <= T168;
    end
    if(T59) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T59) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T120) begin
      pending_ognt_ack <= 1'h1;
    end else if(T103) begin
      pending_ognt_ack <= 1'h1;
    end else if(T211) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T230) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T225) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T238) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T236) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T247) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T245) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T253) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T251) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T59) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T59) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T59) begin
      iacq_data_valid <= T331;
    end else if(T229) begin
      iacq_data_valid <= T325;
    end
    pending_probes <= T425;
  end
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_addr_beat,
    input [1:0] io_in_7_bits_client_xact_id,
    input [3:0] io_in_7_bits_manager_xact_id,
    input  io_in_7_bits_is_builtin_type,
    input [3:0] io_in_7_bits_g_type,
    input [127:0] io_in_7_bits_data,
    input [1:0] io_in_7_bits_client_id,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_addr_beat,
    input [1:0] io_in_6_bits_client_xact_id,
    input [3:0] io_in_6_bits_manager_xact_id,
    input  io_in_6_bits_is_builtin_type,
    input [3:0] io_in_6_bits_g_type,
    input [127:0] io_in_6_bits_data,
    input [1:0] io_in_6_bits_client_id,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_addr_beat,
    input [1:0] io_in_5_bits_client_xact_id,
    input [3:0] io_in_5_bits_manager_xact_id,
    input  io_in_5_bits_is_builtin_type,
    input [3:0] io_in_5_bits_g_type,
    input [127:0] io_in_5_bits_data,
    input [1:0] io_in_5_bits_client_id,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_addr_beat,
    input [1:0] io_in_4_bits_client_xact_id,
    input [3:0] io_in_4_bits_manager_xact_id,
    input  io_in_4_bits_is_builtin_type,
    input [3:0] io_in_4_bits_g_type,
    input [127:0] io_in_4_bits_data,
    input [1:0] io_in_4_bits_client_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_addr_beat,
    input [1:0] io_in_3_bits_client_xact_id,
    input [3:0] io_in_3_bits_manager_xact_id,
    input  io_in_3_bits_is_builtin_type,
    input [3:0] io_in_3_bits_g_type,
    input [127:0] io_in_3_bits_data,
    input [1:0] io_in_3_bits_client_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_addr_beat,
    input [1:0] io_in_2_bits_client_xact_id,
    input [3:0] io_in_2_bits_manager_xact_id,
    input  io_in_2_bits_is_builtin_type,
    input [3:0] io_in_2_bits_g_type,
    input [127:0] io_in_2_bits_data,
    input [1:0] io_in_2_bits_client_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [1:0] io_in_1_bits_client_xact_id,
    input [3:0] io_in_1_bits_manager_xact_id,
    input  io_in_1_bits_is_builtin_type,
    input [3:0] io_in_1_bits_g_type,
    input [127:0] io_in_1_bits_data,
    input [1:0] io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [1:0] io_in_0_bits_client_xact_id,
    input [3:0] io_in_0_bits_manager_xact_id,
    input  io_in_0_bits_is_builtin_type,
    input [3:0] io_in_0_bits_g_type,
    input [127:0] io_in_0_bits_data,
    input [1:0] io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[1:0] io_out_bits_client_xact_id,
    output[3:0] io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[127:0] io_out_bits_data,
    output[1:0] io_out_bits_client_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg [2:0] last_grant;
  wire[2:0] T357;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg [2:0] lockIdx;
  wire[2:0] T358;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  reg  locked;
  wire T359;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  reg [1:0] R59;
  wire[1:0] T360;
  wire[1:0] T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire[1:0] T63;
  wire T64;
  wire[2:0] T65;
  wire[1:0] T66;
  wire T67;
  wire T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[127:0] T76;
  wire[127:0] T77;
  wire[127:0] T78;
  wire T79;
  wire[127:0] T80;
  wire T81;
  wire T82;
  wire[127:0] T83;
  wire[127:0] T84;
  wire T85;
  wire[127:0] T86;
  wire T87;
  wire T88;
  wire T89;
  wire[3:0] T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire T93;
  wire[3:0] T94;
  wire T95;
  wire T96;
  wire[3:0] T97;
  wire[3:0] T98;
  wire T99;
  wire[3:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire[3:0] T118;
  wire[3:0] T119;
  wire[3:0] T120;
  wire T121;
  wire[3:0] T122;
  wire T123;
  wire T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire T127;
  wire[3:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire T135;
  wire[1:0] T136;
  wire T137;
  wire T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[1:0] T146;
  wire[1:0] T147;
  wire[1:0] T148;
  wire T149;
  wire[1:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire T155;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R59 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T28 ? 3'h1 : T1;
  assign T1 = T26 ? 3'h2 : T2;
  assign T2 = T24 ? 3'h3 : T3;
  assign T3 = T22 ? 3'h4 : T4;
  assign T4 = T20 ? 3'h5 : T5;
  assign T5 = T18 ? 3'h6 : T6;
  assign T6 = T14 ? 3'h7 : T7;
  assign T7 = io_in_0_valid ? 3'h0 : T8;
  assign T8 = io_in_1_valid ? 3'h1 : T9;
  assign T9 = io_in_2_valid ? 3'h2 : T10;
  assign T10 = io_in_3_valid ? 3'h3 : T11;
  assign T11 = io_in_4_valid ? 3'h4 : T12;
  assign T12 = io_in_5_valid ? 3'h5 : T13;
  assign T13 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T14 = io_in_7_valid & T15;
  assign T15 = last_grant < 3'h7;
  assign T357 = reset ? 3'h0 : T16;
  assign T16 = T17 ? chosen : last_grant;
  assign T17 = io_out_ready & io_out_valid;
  assign T18 = io_in_6_valid & T19;
  assign T19 = last_grant < 3'h6;
  assign T20 = io_in_5_valid & T21;
  assign T21 = last_grant < 3'h5;
  assign T22 = io_in_4_valid & T23;
  assign T23 = last_grant < 3'h4;
  assign T24 = io_in_3_valid & T25;
  assign T25 = last_grant < 3'h3;
  assign T26 = io_in_2_valid & T27;
  assign T27 = last_grant < 3'h2;
  assign T28 = io_in_1_valid & T29;
  assign T29 = last_grant < 3'h1;
  assign T358 = reset ? 3'h7 : T30;
  assign T30 = T45 ? T31 : lockIdx;
  assign T31 = T44 ? 3'h0 : T32;
  assign T32 = T43 ? 3'h1 : T33;
  assign T33 = T42 ? 3'h2 : T34;
  assign T34 = T41 ? 3'h3 : T35;
  assign T35 = T40 ? 3'h4 : T36;
  assign T36 = T39 ? 3'h5 : T37;
  assign T37 = T38 ? 3'h6 : 3'h7;
  assign T38 = io_in_6_ready & io_in_6_valid;
  assign T39 = io_in_5_ready & io_in_5_valid;
  assign T40 = io_in_4_ready & io_in_4_valid;
  assign T41 = io_in_3_ready & io_in_3_valid;
  assign T42 = io_in_2_ready & io_in_2_valid;
  assign T43 = io_in_1_ready & io_in_1_valid;
  assign T44 = io_in_0_ready & io_in_0_valid;
  assign T45 = T47 & T46;
  assign T46 = locked ^ 1'h1;
  assign T47 = T53 & T48;
  assign T48 = io_out_bits_is_builtin_type ? T52 : T49;
  assign T49 = T51 | T50;
  assign T50 = 4'h1 == io_out_bits_g_type;
  assign T51 = 4'h0 == io_out_bits_g_type;
  assign T52 = 4'h5 == io_out_bits_g_type;
  assign T53 = io_out_ready & io_out_valid;
  assign T359 = reset ? 1'h0 : T54;
  assign T54 = T56 ? 1'h0 : T55;
  assign T55 = T45 ? 1'h1 : locked;
  assign T56 = T53 & T57;
  assign T57 = T58 == 2'h0;
  assign T58 = R59 + 2'h1;
  assign T360 = reset ? 2'h0 : T60;
  assign T60 = T47 ? T58 : R59;
  assign io_out_bits_client_id = T61;
  assign T61 = T75 ? T69 : T62;
  assign T62 = T68 ? T66 : T63;
  assign T63 = T64 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T64 = T65[1'h0:1'h0];
  assign T65 = chosen;
  assign T66 = T67 ? io_in_3_bits_client_id : io_in_2_bits_client_id;
  assign T67 = T65[1'h0:1'h0];
  assign T68 = T65[1'h1:1'h1];
  assign T69 = T74 ? T72 : T70;
  assign T70 = T71 ? io_in_5_bits_client_id : io_in_4_bits_client_id;
  assign T71 = T65[1'h0:1'h0];
  assign T72 = T73 ? io_in_7_bits_client_id : io_in_6_bits_client_id;
  assign T73 = T65[1'h0:1'h0];
  assign T74 = T65[1'h1:1'h1];
  assign T75 = T65[2'h2:2'h2];
  assign io_out_bits_data = T76;
  assign T76 = T89 ? T83 : T77;
  assign T77 = T82 ? T80 : T78;
  assign T78 = T79 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T79 = T65[1'h0:1'h0];
  assign T80 = T81 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T81 = T65[1'h0:1'h0];
  assign T82 = T65[1'h1:1'h1];
  assign T83 = T88 ? T86 : T84;
  assign T84 = T85 ? io_in_5_bits_data : io_in_4_bits_data;
  assign T85 = T65[1'h0:1'h0];
  assign T86 = T87 ? io_in_7_bits_data : io_in_6_bits_data;
  assign T87 = T65[1'h0:1'h0];
  assign T88 = T65[1'h1:1'h1];
  assign T89 = T65[2'h2:2'h2];
  assign io_out_bits_g_type = T90;
  assign T90 = T103 ? T97 : T91;
  assign T91 = T96 ? T94 : T92;
  assign T92 = T93 ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign T93 = T65[1'h0:1'h0];
  assign T94 = T95 ? io_in_3_bits_g_type : io_in_2_bits_g_type;
  assign T95 = T65[1'h0:1'h0];
  assign T96 = T65[1'h1:1'h1];
  assign T97 = T102 ? T100 : T98;
  assign T98 = T99 ? io_in_5_bits_g_type : io_in_4_bits_g_type;
  assign T99 = T65[1'h0:1'h0];
  assign T100 = T101 ? io_in_7_bits_g_type : io_in_6_bits_g_type;
  assign T101 = T65[1'h0:1'h0];
  assign T102 = T65[1'h1:1'h1];
  assign T103 = T65[2'h2:2'h2];
  assign io_out_bits_is_builtin_type = T104;
  assign T104 = T117 ? T111 : T105;
  assign T105 = T110 ? T108 : T106;
  assign T106 = T107 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T107 = T65[1'h0:1'h0];
  assign T108 = T109 ? io_in_3_bits_is_builtin_type : io_in_2_bits_is_builtin_type;
  assign T109 = T65[1'h0:1'h0];
  assign T110 = T65[1'h1:1'h1];
  assign T111 = T116 ? T114 : T112;
  assign T112 = T113 ? io_in_5_bits_is_builtin_type : io_in_4_bits_is_builtin_type;
  assign T113 = T65[1'h0:1'h0];
  assign T114 = T115 ? io_in_7_bits_is_builtin_type : io_in_6_bits_is_builtin_type;
  assign T115 = T65[1'h0:1'h0];
  assign T116 = T65[1'h1:1'h1];
  assign T117 = T65[2'h2:2'h2];
  assign io_out_bits_manager_xact_id = T118;
  assign T118 = T131 ? T125 : T119;
  assign T119 = T124 ? T122 : T120;
  assign T120 = T121 ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign T121 = T65[1'h0:1'h0];
  assign T122 = T123 ? io_in_3_bits_manager_xact_id : io_in_2_bits_manager_xact_id;
  assign T123 = T65[1'h0:1'h0];
  assign T124 = T65[1'h1:1'h1];
  assign T125 = T130 ? T128 : T126;
  assign T126 = T127 ? io_in_5_bits_manager_xact_id : io_in_4_bits_manager_xact_id;
  assign T127 = T65[1'h0:1'h0];
  assign T128 = T129 ? io_in_7_bits_manager_xact_id : io_in_6_bits_manager_xact_id;
  assign T129 = T65[1'h0:1'h0];
  assign T130 = T65[1'h1:1'h1];
  assign T131 = T65[2'h2:2'h2];
  assign io_out_bits_client_xact_id = T132;
  assign T132 = T145 ? T139 : T133;
  assign T133 = T138 ? T136 : T134;
  assign T134 = T135 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T135 = T65[1'h0:1'h0];
  assign T136 = T137 ? io_in_3_bits_client_xact_id : io_in_2_bits_client_xact_id;
  assign T137 = T65[1'h0:1'h0];
  assign T138 = T65[1'h1:1'h1];
  assign T139 = T144 ? T142 : T140;
  assign T140 = T141 ? io_in_5_bits_client_xact_id : io_in_4_bits_client_xact_id;
  assign T141 = T65[1'h0:1'h0];
  assign T142 = T143 ? io_in_7_bits_client_xact_id : io_in_6_bits_client_xact_id;
  assign T143 = T65[1'h0:1'h0];
  assign T144 = T65[1'h1:1'h1];
  assign T145 = T65[2'h2:2'h2];
  assign io_out_bits_addr_beat = T146;
  assign T146 = T159 ? T153 : T147;
  assign T147 = T152 ? T150 : T148;
  assign T148 = T149 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T149 = T65[1'h0:1'h0];
  assign T150 = T151 ? io_in_3_bits_addr_beat : io_in_2_bits_addr_beat;
  assign T151 = T65[1'h0:1'h0];
  assign T152 = T65[1'h1:1'h1];
  assign T153 = T158 ? T156 : T154;
  assign T154 = T155 ? io_in_5_bits_addr_beat : io_in_4_bits_addr_beat;
  assign T155 = T65[1'h0:1'h0];
  assign T156 = T157 ? io_in_7_bits_addr_beat : io_in_6_bits_addr_beat;
  assign T157 = T65[1'h0:1'h0];
  assign T158 = T65[1'h1:1'h1];
  assign T159 = T65[2'h2:2'h2];
  assign io_out_valid = T160;
  assign T160 = T173 ? T167 : T161;
  assign T161 = T166 ? T164 : T162;
  assign T162 = T163 ? io_in_1_valid : io_in_0_valid;
  assign T163 = T65[1'h0:1'h0];
  assign T164 = T165 ? io_in_3_valid : io_in_2_valid;
  assign T165 = T65[1'h0:1'h0];
  assign T166 = T65[1'h1:1'h1];
  assign T167 = T172 ? T170 : T168;
  assign T168 = T169 ? io_in_5_valid : io_in_4_valid;
  assign T169 = T65[1'h0:1'h0];
  assign T170 = T171 ? io_in_7_valid : io_in_6_valid;
  assign T171 = T65[1'h0:1'h0];
  assign T172 = T65[1'h1:1'h1];
  assign T173 = T65[2'h2:2'h2];
  assign io_in_0_ready = T174;
  assign T174 = T175 & io_out_ready;
  assign T175 = locked ? T202 : T176;
  assign T176 = T201 | T177;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T181 | T179;
  assign T179 = io_in_7_valid & T180;
  assign T180 = last_grant < 3'h7;
  assign T181 = T184 | T182;
  assign T182 = io_in_6_valid & T183;
  assign T183 = last_grant < 3'h6;
  assign T184 = T187 | T185;
  assign T185 = io_in_5_valid & T186;
  assign T186 = last_grant < 3'h5;
  assign T187 = T190 | T188;
  assign T188 = io_in_4_valid & T189;
  assign T189 = last_grant < 3'h4;
  assign T190 = T193 | T191;
  assign T191 = io_in_3_valid & T192;
  assign T192 = last_grant < 3'h3;
  assign T193 = T196 | T194;
  assign T194 = io_in_2_valid & T195;
  assign T195 = last_grant < 3'h2;
  assign T196 = T199 | T197;
  assign T197 = io_in_1_valid & T198;
  assign T198 = last_grant < 3'h1;
  assign T199 = io_in_0_valid & T200;
  assign T200 = last_grant < 3'h0;
  assign T201 = last_grant < 3'h0;
  assign T202 = lockIdx == 3'h0;
  assign io_in_1_ready = T203;
  assign T203 = T204 & io_out_ready;
  assign T204 = locked ? T218 : T205;
  assign T205 = T215 | T206;
  assign T206 = T207 ^ 1'h1;
  assign T207 = T208 | io_in_0_valid;
  assign T208 = T209 | T179;
  assign T209 = T210 | T182;
  assign T210 = T211 | T185;
  assign T211 = T212 | T188;
  assign T212 = T213 | T191;
  assign T213 = T214 | T194;
  assign T214 = T199 | T197;
  assign T215 = T217 & T216;
  assign T216 = last_grant < 3'h1;
  assign T217 = T199 ^ 1'h1;
  assign T218 = lockIdx == 3'h1;
  assign io_in_2_ready = T219;
  assign T219 = T220 & io_out_ready;
  assign T220 = locked ? T236 : T221;
  assign T221 = T232 | T222;
  assign T222 = T223 ^ 1'h1;
  assign T223 = T224 | io_in_1_valid;
  assign T224 = T225 | io_in_0_valid;
  assign T225 = T226 | T179;
  assign T226 = T227 | T182;
  assign T227 = T228 | T185;
  assign T228 = T229 | T188;
  assign T229 = T230 | T191;
  assign T230 = T231 | T194;
  assign T231 = T199 | T197;
  assign T232 = T234 & T233;
  assign T233 = last_grant < 3'h2;
  assign T234 = T235 ^ 1'h1;
  assign T235 = T199 | T197;
  assign T236 = lockIdx == 3'h2;
  assign io_in_3_ready = T237;
  assign T237 = T238 & io_out_ready;
  assign T238 = locked ? T256 : T239;
  assign T239 = T251 | T240;
  assign T240 = T241 ^ 1'h1;
  assign T241 = T242 | io_in_2_valid;
  assign T242 = T243 | io_in_1_valid;
  assign T243 = T244 | io_in_0_valid;
  assign T244 = T245 | T179;
  assign T245 = T246 | T182;
  assign T246 = T247 | T185;
  assign T247 = T248 | T188;
  assign T248 = T249 | T191;
  assign T249 = T250 | T194;
  assign T250 = T199 | T197;
  assign T251 = T253 & T252;
  assign T252 = last_grant < 3'h3;
  assign T253 = T254 ^ 1'h1;
  assign T254 = T255 | T194;
  assign T255 = T199 | T197;
  assign T256 = lockIdx == 3'h3;
  assign io_in_4_ready = T257;
  assign T257 = T258 & io_out_ready;
  assign T258 = locked ? T278 : T259;
  assign T259 = T272 | T260;
  assign T260 = T261 ^ 1'h1;
  assign T261 = T262 | io_in_3_valid;
  assign T262 = T263 | io_in_2_valid;
  assign T263 = T264 | io_in_1_valid;
  assign T264 = T265 | io_in_0_valid;
  assign T265 = T266 | T179;
  assign T266 = T267 | T182;
  assign T267 = T268 | T185;
  assign T268 = T269 | T188;
  assign T269 = T270 | T191;
  assign T270 = T271 | T194;
  assign T271 = T199 | T197;
  assign T272 = T274 & T273;
  assign T273 = last_grant < 3'h4;
  assign T274 = T275 ^ 1'h1;
  assign T275 = T276 | T191;
  assign T276 = T277 | T194;
  assign T277 = T199 | T197;
  assign T278 = lockIdx == 3'h4;
  assign io_in_5_ready = T279;
  assign T279 = T280 & io_out_ready;
  assign T280 = locked ? T302 : T281;
  assign T281 = T295 | T282;
  assign T282 = T283 ^ 1'h1;
  assign T283 = T284 | io_in_4_valid;
  assign T284 = T285 | io_in_3_valid;
  assign T285 = T286 | io_in_2_valid;
  assign T286 = T287 | io_in_1_valid;
  assign T287 = T288 | io_in_0_valid;
  assign T288 = T289 | T179;
  assign T289 = T290 | T182;
  assign T290 = T291 | T185;
  assign T291 = T292 | T188;
  assign T292 = T293 | T191;
  assign T293 = T294 | T194;
  assign T294 = T199 | T197;
  assign T295 = T297 & T296;
  assign T296 = last_grant < 3'h5;
  assign T297 = T298 ^ 1'h1;
  assign T298 = T299 | T188;
  assign T299 = T300 | T191;
  assign T300 = T301 | T194;
  assign T301 = T199 | T197;
  assign T302 = lockIdx == 3'h5;
  assign io_in_6_ready = T303;
  assign T303 = T304 & io_out_ready;
  assign T304 = locked ? T328 : T305;
  assign T305 = T320 | T306;
  assign T306 = T307 ^ 1'h1;
  assign T307 = T308 | io_in_5_valid;
  assign T308 = T309 | io_in_4_valid;
  assign T309 = T310 | io_in_3_valid;
  assign T310 = T311 | io_in_2_valid;
  assign T311 = T312 | io_in_1_valid;
  assign T312 = T313 | io_in_0_valid;
  assign T313 = T314 | T179;
  assign T314 = T315 | T182;
  assign T315 = T316 | T185;
  assign T316 = T317 | T188;
  assign T317 = T318 | T191;
  assign T318 = T319 | T194;
  assign T319 = T199 | T197;
  assign T320 = T322 & T321;
  assign T321 = last_grant < 3'h6;
  assign T322 = T323 ^ 1'h1;
  assign T323 = T324 | T185;
  assign T324 = T325 | T188;
  assign T325 = T326 | T191;
  assign T326 = T327 | T194;
  assign T327 = T199 | T197;
  assign T328 = lockIdx == 3'h6;
  assign io_in_7_ready = T329;
  assign T329 = T330 & io_out_ready;
  assign T330 = locked ? T356 : T331;
  assign T331 = T347 | T332;
  assign T332 = T333 ^ 1'h1;
  assign T333 = T334 | io_in_6_valid;
  assign T334 = T335 | io_in_5_valid;
  assign T335 = T336 | io_in_4_valid;
  assign T336 = T337 | io_in_3_valid;
  assign T337 = T338 | io_in_2_valid;
  assign T338 = T339 | io_in_1_valid;
  assign T339 = T340 | io_in_0_valid;
  assign T340 = T341 | T179;
  assign T341 = T342 | T182;
  assign T342 = T343 | T185;
  assign T343 = T344 | T188;
  assign T344 = T345 | T191;
  assign T345 = T346 | T194;
  assign T346 = T199 | T197;
  assign T347 = T349 & T348;
  assign T348 = last_grant < 3'h7;
  assign T349 = T350 ^ 1'h1;
  assign T350 = T351 | T182;
  assign T351 = T352 | T185;
  assign T352 = T353 | T188;
  assign T353 = T354 | T191;
  assign T354 = T355 | T194;
  assign T355 = T199 | T197;
  assign T356 = lockIdx == 3'h7;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T17) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h7;
    end else if(T45) begin
      lockIdx <= T31;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T56) begin
      locked <= 1'h0;
    end else if(T45) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R59 <= 2'h0;
    end else if(T47) begin
      R59 <= T58;
    end
  end
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [25:0] io_in_7_bits_addr_block,
    input [1:0] io_in_7_bits_p_type,
    input [1:0] io_in_7_bits_client_id,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [25:0] io_in_6_bits_addr_block,
    input [1:0] io_in_6_bits_p_type,
    input [1:0] io_in_6_bits_client_id,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [25:0] io_in_5_bits_addr_block,
    input [1:0] io_in_5_bits_p_type,
    input [1:0] io_in_5_bits_client_id,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [25:0] io_in_4_bits_addr_block,
    input [1:0] io_in_4_bits_p_type,
    input [1:0] io_in_4_bits_client_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [25:0] io_in_3_bits_addr_block,
    input [1:0] io_in_3_bits_p_type,
    input [1:0] io_in_3_bits_client_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [1:0] io_in_2_bits_p_type,
    input [1:0] io_in_2_bits_client_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_p_type,
    input [1:0] io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_p_type,
    input [1:0] io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_p_type,
    output[1:0] io_out_bits_client_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg [2:0] last_grant;
  wire[2:0] T276;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg [2:0] lockIdx;
  wire[2:0] T277;
  reg  locked;
  wire T278;
  wire T30;
  wire T31;
  wire T32;
  wire[1:0] T33;
  reg [1:0] R34;
  wire[1:0] T279;
  wire T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire[2:0] T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[25:0] T65;
  wire[25:0] T66;
  wire[25:0] T67;
  wire T68;
  wire[25:0] T69;
  wire T70;
  wire T71;
  wire[25:0] T72;
  wire[25:0] T73;
  wire T74;
  wire[25:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R34 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T28 ? 3'h1 : T1;
  assign T1 = T26 ? 3'h2 : T2;
  assign T2 = T24 ? 3'h3 : T3;
  assign T3 = T22 ? 3'h4 : T4;
  assign T4 = T20 ? 3'h5 : T5;
  assign T5 = T18 ? 3'h6 : T6;
  assign T6 = T14 ? 3'h7 : T7;
  assign T7 = io_in_0_valid ? 3'h0 : T8;
  assign T8 = io_in_1_valid ? 3'h1 : T9;
  assign T9 = io_in_2_valid ? 3'h2 : T10;
  assign T10 = io_in_3_valid ? 3'h3 : T11;
  assign T11 = io_in_4_valid ? 3'h4 : T12;
  assign T12 = io_in_5_valid ? 3'h5 : T13;
  assign T13 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T14 = io_in_7_valid & T15;
  assign T15 = last_grant < 3'h7;
  assign T276 = reset ? 3'h0 : T16;
  assign T16 = T17 ? chosen : last_grant;
  assign T17 = io_out_ready & io_out_valid;
  assign T18 = io_in_6_valid & T19;
  assign T19 = last_grant < 3'h6;
  assign T20 = io_in_5_valid & T21;
  assign T21 = last_grant < 3'h5;
  assign T22 = io_in_4_valid & T23;
  assign T23 = last_grant < 3'h4;
  assign T24 = io_in_3_valid & T25;
  assign T25 = last_grant < 3'h3;
  assign T26 = io_in_2_valid & T27;
  assign T27 = last_grant < 3'h2;
  assign T28 = io_in_1_valid & T29;
  assign T29 = last_grant < 3'h1;
  assign T277 = reset ? 3'h7 : lockIdx;
  assign T278 = reset ? 1'h0 : T30;
  assign T30 = T31 ? 1'h0 : locked;
  assign T31 = T35 & T32;
  assign T32 = T33 == 2'h0;
  assign T33 = R34 + 2'h1;
  assign T279 = reset ? 2'h0 : R34;
  assign T35 = io_out_ready & io_out_valid;
  assign io_out_bits_client_id = T36;
  assign T36 = T50 ? T44 : T37;
  assign T37 = T43 ? T41 : T38;
  assign T38 = T39 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T39 = T40[1'h0:1'h0];
  assign T40 = chosen;
  assign T41 = T42 ? io_in_3_bits_client_id : io_in_2_bits_client_id;
  assign T42 = T40[1'h0:1'h0];
  assign T43 = T40[1'h1:1'h1];
  assign T44 = T49 ? T47 : T45;
  assign T45 = T46 ? io_in_5_bits_client_id : io_in_4_bits_client_id;
  assign T46 = T40[1'h0:1'h0];
  assign T47 = T48 ? io_in_7_bits_client_id : io_in_6_bits_client_id;
  assign T48 = T40[1'h0:1'h0];
  assign T49 = T40[1'h1:1'h1];
  assign T50 = T40[2'h2:2'h2];
  assign io_out_bits_p_type = T51;
  assign T51 = T64 ? T58 : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_p_type : io_in_0_bits_p_type;
  assign T54 = T40[1'h0:1'h0];
  assign T55 = T56 ? io_in_3_bits_p_type : io_in_2_bits_p_type;
  assign T56 = T40[1'h0:1'h0];
  assign T57 = T40[1'h1:1'h1];
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_5_bits_p_type : io_in_4_bits_p_type;
  assign T60 = T40[1'h0:1'h0];
  assign T61 = T62 ? io_in_7_bits_p_type : io_in_6_bits_p_type;
  assign T62 = T40[1'h0:1'h0];
  assign T63 = T40[1'h1:1'h1];
  assign T64 = T40[2'h2:2'h2];
  assign io_out_bits_addr_block = T65;
  assign T65 = T78 ? T72 : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T68 = T40[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_addr_block : io_in_2_bits_addr_block;
  assign T70 = T40[1'h0:1'h0];
  assign T71 = T40[1'h1:1'h1];
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74 ? io_in_5_bits_addr_block : io_in_4_bits_addr_block;
  assign T74 = T40[1'h0:1'h0];
  assign T75 = T76 ? io_in_7_bits_addr_block : io_in_6_bits_addr_block;
  assign T76 = T40[1'h0:1'h0];
  assign T77 = T40[1'h1:1'h1];
  assign T78 = T40[2'h2:2'h2];
  assign io_out_valid = T79;
  assign T79 = T92 ? T86 : T80;
  assign T80 = T85 ? T83 : T81;
  assign T81 = T82 ? io_in_1_valid : io_in_0_valid;
  assign T82 = T40[1'h0:1'h0];
  assign T83 = T84 ? io_in_3_valid : io_in_2_valid;
  assign T84 = T40[1'h0:1'h0];
  assign T85 = T40[1'h1:1'h1];
  assign T86 = T91 ? T89 : T87;
  assign T87 = T88 ? io_in_5_valid : io_in_4_valid;
  assign T88 = T40[1'h0:1'h0];
  assign T89 = T90 ? io_in_7_valid : io_in_6_valid;
  assign T90 = T40[1'h0:1'h0];
  assign T91 = T40[1'h1:1'h1];
  assign T92 = T40[2'h2:2'h2];
  assign io_in_0_ready = T93;
  assign T93 = T94 & io_out_ready;
  assign T94 = locked ? T121 : T95;
  assign T95 = T120 | T96;
  assign T96 = T97 ^ 1'h1;
  assign T97 = T100 | T98;
  assign T98 = io_in_7_valid & T99;
  assign T99 = last_grant < 3'h7;
  assign T100 = T103 | T101;
  assign T101 = io_in_6_valid & T102;
  assign T102 = last_grant < 3'h6;
  assign T103 = T106 | T104;
  assign T104 = io_in_5_valid & T105;
  assign T105 = last_grant < 3'h5;
  assign T106 = T109 | T107;
  assign T107 = io_in_4_valid & T108;
  assign T108 = last_grant < 3'h4;
  assign T109 = T112 | T110;
  assign T110 = io_in_3_valid & T111;
  assign T111 = last_grant < 3'h3;
  assign T112 = T115 | T113;
  assign T113 = io_in_2_valid & T114;
  assign T114 = last_grant < 3'h2;
  assign T115 = T118 | T116;
  assign T116 = io_in_1_valid & T117;
  assign T117 = last_grant < 3'h1;
  assign T118 = io_in_0_valid & T119;
  assign T119 = last_grant < 3'h0;
  assign T120 = last_grant < 3'h0;
  assign T121 = lockIdx == 3'h0;
  assign io_in_1_ready = T122;
  assign T122 = T123 & io_out_ready;
  assign T123 = locked ? T137 : T124;
  assign T124 = T134 | T125;
  assign T125 = T126 ^ 1'h1;
  assign T126 = T127 | io_in_0_valid;
  assign T127 = T128 | T98;
  assign T128 = T129 | T101;
  assign T129 = T130 | T104;
  assign T130 = T131 | T107;
  assign T131 = T132 | T110;
  assign T132 = T133 | T113;
  assign T133 = T118 | T116;
  assign T134 = T136 & T135;
  assign T135 = last_grant < 3'h1;
  assign T136 = T118 ^ 1'h1;
  assign T137 = lockIdx == 3'h1;
  assign io_in_2_ready = T138;
  assign T138 = T139 & io_out_ready;
  assign T139 = locked ? T155 : T140;
  assign T140 = T151 | T141;
  assign T141 = T142 ^ 1'h1;
  assign T142 = T143 | io_in_1_valid;
  assign T143 = T144 | io_in_0_valid;
  assign T144 = T145 | T98;
  assign T145 = T146 | T101;
  assign T146 = T147 | T104;
  assign T147 = T148 | T107;
  assign T148 = T149 | T110;
  assign T149 = T150 | T113;
  assign T150 = T118 | T116;
  assign T151 = T153 & T152;
  assign T152 = last_grant < 3'h2;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T118 | T116;
  assign T155 = lockIdx == 3'h2;
  assign io_in_3_ready = T156;
  assign T156 = T157 & io_out_ready;
  assign T157 = locked ? T175 : T158;
  assign T158 = T170 | T159;
  assign T159 = T160 ^ 1'h1;
  assign T160 = T161 | io_in_2_valid;
  assign T161 = T162 | io_in_1_valid;
  assign T162 = T163 | io_in_0_valid;
  assign T163 = T164 | T98;
  assign T164 = T165 | T101;
  assign T165 = T166 | T104;
  assign T166 = T167 | T107;
  assign T167 = T168 | T110;
  assign T168 = T169 | T113;
  assign T169 = T118 | T116;
  assign T170 = T172 & T171;
  assign T171 = last_grant < 3'h3;
  assign T172 = T173 ^ 1'h1;
  assign T173 = T174 | T113;
  assign T174 = T118 | T116;
  assign T175 = lockIdx == 3'h3;
  assign io_in_4_ready = T176;
  assign T176 = T177 & io_out_ready;
  assign T177 = locked ? T197 : T178;
  assign T178 = T191 | T179;
  assign T179 = T180 ^ 1'h1;
  assign T180 = T181 | io_in_3_valid;
  assign T181 = T182 | io_in_2_valid;
  assign T182 = T183 | io_in_1_valid;
  assign T183 = T184 | io_in_0_valid;
  assign T184 = T185 | T98;
  assign T185 = T186 | T101;
  assign T186 = T187 | T104;
  assign T187 = T188 | T107;
  assign T188 = T189 | T110;
  assign T189 = T190 | T113;
  assign T190 = T118 | T116;
  assign T191 = T193 & T192;
  assign T192 = last_grant < 3'h4;
  assign T193 = T194 ^ 1'h1;
  assign T194 = T195 | T110;
  assign T195 = T196 | T113;
  assign T196 = T118 | T116;
  assign T197 = lockIdx == 3'h4;
  assign io_in_5_ready = T198;
  assign T198 = T199 & io_out_ready;
  assign T199 = locked ? T221 : T200;
  assign T200 = T214 | T201;
  assign T201 = T202 ^ 1'h1;
  assign T202 = T203 | io_in_4_valid;
  assign T203 = T204 | io_in_3_valid;
  assign T204 = T205 | io_in_2_valid;
  assign T205 = T206 | io_in_1_valid;
  assign T206 = T207 | io_in_0_valid;
  assign T207 = T208 | T98;
  assign T208 = T209 | T101;
  assign T209 = T210 | T104;
  assign T210 = T211 | T107;
  assign T211 = T212 | T110;
  assign T212 = T213 | T113;
  assign T213 = T118 | T116;
  assign T214 = T216 & T215;
  assign T215 = last_grant < 3'h5;
  assign T216 = T217 ^ 1'h1;
  assign T217 = T218 | T107;
  assign T218 = T219 | T110;
  assign T219 = T220 | T113;
  assign T220 = T118 | T116;
  assign T221 = lockIdx == 3'h5;
  assign io_in_6_ready = T222;
  assign T222 = T223 & io_out_ready;
  assign T223 = locked ? T247 : T224;
  assign T224 = T239 | T225;
  assign T225 = T226 ^ 1'h1;
  assign T226 = T227 | io_in_5_valid;
  assign T227 = T228 | io_in_4_valid;
  assign T228 = T229 | io_in_3_valid;
  assign T229 = T230 | io_in_2_valid;
  assign T230 = T231 | io_in_1_valid;
  assign T231 = T232 | io_in_0_valid;
  assign T232 = T233 | T98;
  assign T233 = T234 | T101;
  assign T234 = T235 | T104;
  assign T235 = T236 | T107;
  assign T236 = T237 | T110;
  assign T237 = T238 | T113;
  assign T238 = T118 | T116;
  assign T239 = T241 & T240;
  assign T240 = last_grant < 3'h6;
  assign T241 = T242 ^ 1'h1;
  assign T242 = T243 | T104;
  assign T243 = T244 | T107;
  assign T244 = T245 | T110;
  assign T245 = T246 | T113;
  assign T246 = T118 | T116;
  assign T247 = lockIdx == 3'h6;
  assign io_in_7_ready = T248;
  assign T248 = T249 & io_out_ready;
  assign T249 = locked ? T275 : T250;
  assign T250 = T266 | T251;
  assign T251 = T252 ^ 1'h1;
  assign T252 = T253 | io_in_6_valid;
  assign T253 = T254 | io_in_5_valid;
  assign T254 = T255 | io_in_4_valid;
  assign T255 = T256 | io_in_3_valid;
  assign T256 = T257 | io_in_2_valid;
  assign T257 = T258 | io_in_1_valid;
  assign T258 = T259 | io_in_0_valid;
  assign T259 = T260 | T98;
  assign T260 = T261 | T101;
  assign T261 = T262 | T104;
  assign T262 = T263 | T107;
  assign T263 = T264 | T110;
  assign T264 = T265 | T113;
  assign T265 = T118 | T116;
  assign T266 = T268 & T267;
  assign T267 = last_grant < 3'h7;
  assign T268 = T269 ^ 1'h1;
  assign T269 = T270 | T101;
  assign T270 = T271 | T104;
  assign T271 = T272 | T107;
  assign T272 = T273 | T110;
  assign T273 = T274 | T113;
  assign T274 = T118 | T116;
  assign T275 = lockIdx == 3'h7;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T17) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h7;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T31) begin
      locked <= 1'h0;
    end
    if(reset) begin
      R34 <= 2'h0;
    end
  end
endmodule

module LockingRRArbiter_5(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [25:0] io_in_7_bits_addr_block,
    input [3:0] io_in_7_bits_client_xact_id,
    input [1:0] io_in_7_bits_addr_beat,
    input  io_in_7_bits_is_builtin_type,
    input [2:0] io_in_7_bits_a_type,
    input [16:0] io_in_7_bits_union,
    input [3:0] io_in_7_bits_data,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [25:0] io_in_6_bits_addr_block,
    input [3:0] io_in_6_bits_client_xact_id,
    input [1:0] io_in_6_bits_addr_beat,
    input  io_in_6_bits_is_builtin_type,
    input [2:0] io_in_6_bits_a_type,
    input [16:0] io_in_6_bits_union,
    input [3:0] io_in_6_bits_data,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [25:0] io_in_5_bits_addr_block,
    input [3:0] io_in_5_bits_client_xact_id,
    input [1:0] io_in_5_bits_addr_beat,
    input  io_in_5_bits_is_builtin_type,
    input [2:0] io_in_5_bits_a_type,
    input [16:0] io_in_5_bits_union,
    input [3:0] io_in_5_bits_data,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [25:0] io_in_4_bits_addr_block,
    input [3:0] io_in_4_bits_client_xact_id,
    input [1:0] io_in_4_bits_addr_beat,
    input  io_in_4_bits_is_builtin_type,
    input [2:0] io_in_4_bits_a_type,
    input [16:0] io_in_4_bits_union,
    input [3:0] io_in_4_bits_data,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [25:0] io_in_3_bits_addr_block,
    input [3:0] io_in_3_bits_client_xact_id,
    input [1:0] io_in_3_bits_addr_beat,
    input  io_in_3_bits_is_builtin_type,
    input [2:0] io_in_3_bits_a_type,
    input [16:0] io_in_3_bits_union,
    input [3:0] io_in_3_bits_data,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [3:0] io_in_2_bits_client_xact_id,
    input [1:0] io_in_2_bits_addr_beat,
    input  io_in_2_bits_is_builtin_type,
    input [2:0] io_in_2_bits_a_type,
    input [16:0] io_in_2_bits_union,
    input [3:0] io_in_2_bits_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [3:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [3:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [3:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [3:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[3:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[3:0] io_out_bits_data,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg [2:0] last_grant;
  wire[2:0] T354;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg [2:0] lockIdx;
  wire[2:0] T355;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  reg  locked;
  wire T356;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  reg [1:0] R56;
  wire[1:0] T357;
  wire[1:0] T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T60;
  wire T61;
  wire[2:0] T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire[3:0] T67;
  wire T68;
  wire[3:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire[16:0] T73;
  wire[16:0] T74;
  wire[16:0] T75;
  wire T76;
  wire[16:0] T77;
  wire T78;
  wire T79;
  wire[16:0] T80;
  wire[16:0] T81;
  wire T82;
  wire[16:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire[2:0] T87;
  wire[2:0] T88;
  wire[2:0] T89;
  wire T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire T96;
  wire[2:0] T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire[1:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire[3:0] T129;
  wire[3:0] T130;
  wire[3:0] T131;
  wire T132;
  wire[3:0] T133;
  wire T134;
  wire T135;
  wire[3:0] T136;
  wire[3:0] T137;
  wire T138;
  wire[3:0] T139;
  wire T140;
  wire T141;
  wire T142;
  wire[25:0] T143;
  wire[25:0] T144;
  wire[25:0] T145;
  wire T146;
  wire[25:0] T147;
  wire T148;
  wire T149;
  wire[25:0] T150;
  wire[25:0] T151;
  wire T152;
  wire[25:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R56 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T28 ? 3'h1 : T1;
  assign T1 = T26 ? 3'h2 : T2;
  assign T2 = T24 ? 3'h3 : T3;
  assign T3 = T22 ? 3'h4 : T4;
  assign T4 = T20 ? 3'h5 : T5;
  assign T5 = T18 ? 3'h6 : T6;
  assign T6 = T14 ? 3'h7 : T7;
  assign T7 = io_in_0_valid ? 3'h0 : T8;
  assign T8 = io_in_1_valid ? 3'h1 : T9;
  assign T9 = io_in_2_valid ? 3'h2 : T10;
  assign T10 = io_in_3_valid ? 3'h3 : T11;
  assign T11 = io_in_4_valid ? 3'h4 : T12;
  assign T12 = io_in_5_valid ? 3'h5 : T13;
  assign T13 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T14 = io_in_7_valid & T15;
  assign T15 = last_grant < 3'h7;
  assign T354 = reset ? 3'h0 : T16;
  assign T16 = T17 ? chosen : last_grant;
  assign T17 = io_out_ready & io_out_valid;
  assign T18 = io_in_6_valid & T19;
  assign T19 = last_grant < 3'h6;
  assign T20 = io_in_5_valid & T21;
  assign T21 = last_grant < 3'h5;
  assign T22 = io_in_4_valid & T23;
  assign T23 = last_grant < 3'h4;
  assign T24 = io_in_3_valid & T25;
  assign T25 = last_grant < 3'h3;
  assign T26 = io_in_2_valid & T27;
  assign T27 = last_grant < 3'h2;
  assign T28 = io_in_1_valid & T29;
  assign T29 = last_grant < 3'h1;
  assign T355 = reset ? 3'h7 : T30;
  assign T30 = T45 ? T31 : lockIdx;
  assign T31 = T44 ? 3'h0 : T32;
  assign T32 = T43 ? 3'h1 : T33;
  assign T33 = T42 ? 3'h2 : T34;
  assign T34 = T41 ? 3'h3 : T35;
  assign T35 = T40 ? 3'h4 : T36;
  assign T36 = T39 ? 3'h5 : T37;
  assign T37 = T38 ? 3'h6 : 3'h7;
  assign T38 = io_in_6_ready & io_in_6_valid;
  assign T39 = io_in_5_ready & io_in_5_valid;
  assign T40 = io_in_4_ready & io_in_4_valid;
  assign T41 = io_in_3_ready & io_in_3_valid;
  assign T42 = io_in_2_ready & io_in_2_valid;
  assign T43 = io_in_1_ready & io_in_1_valid;
  assign T44 = io_in_0_ready & io_in_0_valid;
  assign T45 = T47 & T46;
  assign T46 = locked ^ 1'h1;
  assign T47 = T50 & T48;
  assign T48 = io_out_bits_is_builtin_type & T49;
  assign T49 = 3'h3 == io_out_bits_a_type;
  assign T50 = io_out_ready & io_out_valid;
  assign T356 = reset ? 1'h0 : T51;
  assign T51 = T53 ? 1'h0 : T52;
  assign T52 = T45 ? 1'h1 : locked;
  assign T53 = T50 & T54;
  assign T54 = T55 == 2'h0;
  assign T55 = R56 + 2'h1;
  assign T357 = reset ? 2'h0 : T57;
  assign T57 = T47 ? T55 : R56;
  assign io_out_bits_data = T58;
  assign T58 = T72 ? T66 : T59;
  assign T59 = T65 ? T63 : T60;
  assign T60 = T61 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T61 = T62[1'h0:1'h0];
  assign T62 = chosen;
  assign T63 = T64 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T64 = T62[1'h0:1'h0];
  assign T65 = T62[1'h1:1'h1];
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_5_bits_data : io_in_4_bits_data;
  assign T68 = T62[1'h0:1'h0];
  assign T69 = T70 ? io_in_7_bits_data : io_in_6_bits_data;
  assign T70 = T62[1'h0:1'h0];
  assign T71 = T62[1'h1:1'h1];
  assign T72 = T62[2'h2:2'h2];
  assign io_out_bits_union = T73;
  assign T73 = T86 ? T80 : T74;
  assign T74 = T79 ? T77 : T75;
  assign T75 = T76 ? io_in_1_bits_union : io_in_0_bits_union;
  assign T76 = T62[1'h0:1'h0];
  assign T77 = T78 ? io_in_3_bits_union : io_in_2_bits_union;
  assign T78 = T62[1'h0:1'h0];
  assign T79 = T62[1'h1:1'h1];
  assign T80 = T85 ? T83 : T81;
  assign T81 = T82 ? io_in_5_bits_union : io_in_4_bits_union;
  assign T82 = T62[1'h0:1'h0];
  assign T83 = T84 ? io_in_7_bits_union : io_in_6_bits_union;
  assign T84 = T62[1'h0:1'h0];
  assign T85 = T62[1'h1:1'h1];
  assign T86 = T62[2'h2:2'h2];
  assign io_out_bits_a_type = T87;
  assign T87 = T100 ? T94 : T88;
  assign T88 = T93 ? T91 : T89;
  assign T89 = T90 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign T90 = T62[1'h0:1'h0];
  assign T91 = T92 ? io_in_3_bits_a_type : io_in_2_bits_a_type;
  assign T92 = T62[1'h0:1'h0];
  assign T93 = T62[1'h1:1'h1];
  assign T94 = T99 ? T97 : T95;
  assign T95 = T96 ? io_in_5_bits_a_type : io_in_4_bits_a_type;
  assign T96 = T62[1'h0:1'h0];
  assign T97 = T98 ? io_in_7_bits_a_type : io_in_6_bits_a_type;
  assign T98 = T62[1'h0:1'h0];
  assign T99 = T62[1'h1:1'h1];
  assign T100 = T62[2'h2:2'h2];
  assign io_out_bits_is_builtin_type = T101;
  assign T101 = T114 ? T108 : T102;
  assign T102 = T107 ? T105 : T103;
  assign T103 = T104 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T104 = T62[1'h0:1'h0];
  assign T105 = T106 ? io_in_3_bits_is_builtin_type : io_in_2_bits_is_builtin_type;
  assign T106 = T62[1'h0:1'h0];
  assign T107 = T62[1'h1:1'h1];
  assign T108 = T113 ? T111 : T109;
  assign T109 = T110 ? io_in_5_bits_is_builtin_type : io_in_4_bits_is_builtin_type;
  assign T110 = T62[1'h0:1'h0];
  assign T111 = T112 ? io_in_7_bits_is_builtin_type : io_in_6_bits_is_builtin_type;
  assign T112 = T62[1'h0:1'h0];
  assign T113 = T62[1'h1:1'h1];
  assign T114 = T62[2'h2:2'h2];
  assign io_out_bits_addr_beat = T115;
  assign T115 = T128 ? T122 : T116;
  assign T116 = T121 ? T119 : T117;
  assign T117 = T118 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T118 = T62[1'h0:1'h0];
  assign T119 = T120 ? io_in_3_bits_addr_beat : io_in_2_bits_addr_beat;
  assign T120 = T62[1'h0:1'h0];
  assign T121 = T62[1'h1:1'h1];
  assign T122 = T127 ? T125 : T123;
  assign T123 = T124 ? io_in_5_bits_addr_beat : io_in_4_bits_addr_beat;
  assign T124 = T62[1'h0:1'h0];
  assign T125 = T126 ? io_in_7_bits_addr_beat : io_in_6_bits_addr_beat;
  assign T126 = T62[1'h0:1'h0];
  assign T127 = T62[1'h1:1'h1];
  assign T128 = T62[2'h2:2'h2];
  assign io_out_bits_client_xact_id = T129;
  assign T129 = T142 ? T136 : T130;
  assign T130 = T135 ? T133 : T131;
  assign T131 = T132 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T132 = T62[1'h0:1'h0];
  assign T133 = T134 ? io_in_3_bits_client_xact_id : io_in_2_bits_client_xact_id;
  assign T134 = T62[1'h0:1'h0];
  assign T135 = T62[1'h1:1'h1];
  assign T136 = T141 ? T139 : T137;
  assign T137 = T138 ? io_in_5_bits_client_xact_id : io_in_4_bits_client_xact_id;
  assign T138 = T62[1'h0:1'h0];
  assign T139 = T140 ? io_in_7_bits_client_xact_id : io_in_6_bits_client_xact_id;
  assign T140 = T62[1'h0:1'h0];
  assign T141 = T62[1'h1:1'h1];
  assign T142 = T62[2'h2:2'h2];
  assign io_out_bits_addr_block = T143;
  assign T143 = T156 ? T150 : T144;
  assign T144 = T149 ? T147 : T145;
  assign T145 = T146 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T146 = T62[1'h0:1'h0];
  assign T147 = T148 ? io_in_3_bits_addr_block : io_in_2_bits_addr_block;
  assign T148 = T62[1'h0:1'h0];
  assign T149 = T62[1'h1:1'h1];
  assign T150 = T155 ? T153 : T151;
  assign T151 = T152 ? io_in_5_bits_addr_block : io_in_4_bits_addr_block;
  assign T152 = T62[1'h0:1'h0];
  assign T153 = T154 ? io_in_7_bits_addr_block : io_in_6_bits_addr_block;
  assign T154 = T62[1'h0:1'h0];
  assign T155 = T62[1'h1:1'h1];
  assign T156 = T62[2'h2:2'h2];
  assign io_out_valid = T157;
  assign T157 = T170 ? T164 : T158;
  assign T158 = T163 ? T161 : T159;
  assign T159 = T160 ? io_in_1_valid : io_in_0_valid;
  assign T160 = T62[1'h0:1'h0];
  assign T161 = T162 ? io_in_3_valid : io_in_2_valid;
  assign T162 = T62[1'h0:1'h0];
  assign T163 = T62[1'h1:1'h1];
  assign T164 = T169 ? T167 : T165;
  assign T165 = T166 ? io_in_5_valid : io_in_4_valid;
  assign T166 = T62[1'h0:1'h0];
  assign T167 = T168 ? io_in_7_valid : io_in_6_valid;
  assign T168 = T62[1'h0:1'h0];
  assign T169 = T62[1'h1:1'h1];
  assign T170 = T62[2'h2:2'h2];
  assign io_in_0_ready = T171;
  assign T171 = T172 & io_out_ready;
  assign T172 = locked ? T199 : T173;
  assign T173 = T198 | T174;
  assign T174 = T175 ^ 1'h1;
  assign T175 = T178 | T176;
  assign T176 = io_in_7_valid & T177;
  assign T177 = last_grant < 3'h7;
  assign T178 = T181 | T179;
  assign T179 = io_in_6_valid & T180;
  assign T180 = last_grant < 3'h6;
  assign T181 = T184 | T182;
  assign T182 = io_in_5_valid & T183;
  assign T183 = last_grant < 3'h5;
  assign T184 = T187 | T185;
  assign T185 = io_in_4_valid & T186;
  assign T186 = last_grant < 3'h4;
  assign T187 = T190 | T188;
  assign T188 = io_in_3_valid & T189;
  assign T189 = last_grant < 3'h3;
  assign T190 = T193 | T191;
  assign T191 = io_in_2_valid & T192;
  assign T192 = last_grant < 3'h2;
  assign T193 = T196 | T194;
  assign T194 = io_in_1_valid & T195;
  assign T195 = last_grant < 3'h1;
  assign T196 = io_in_0_valid & T197;
  assign T197 = last_grant < 3'h0;
  assign T198 = last_grant < 3'h0;
  assign T199 = lockIdx == 3'h0;
  assign io_in_1_ready = T200;
  assign T200 = T201 & io_out_ready;
  assign T201 = locked ? T215 : T202;
  assign T202 = T212 | T203;
  assign T203 = T204 ^ 1'h1;
  assign T204 = T205 | io_in_0_valid;
  assign T205 = T206 | T176;
  assign T206 = T207 | T179;
  assign T207 = T208 | T182;
  assign T208 = T209 | T185;
  assign T209 = T210 | T188;
  assign T210 = T211 | T191;
  assign T211 = T196 | T194;
  assign T212 = T214 & T213;
  assign T213 = last_grant < 3'h1;
  assign T214 = T196 ^ 1'h1;
  assign T215 = lockIdx == 3'h1;
  assign io_in_2_ready = T216;
  assign T216 = T217 & io_out_ready;
  assign T217 = locked ? T233 : T218;
  assign T218 = T229 | T219;
  assign T219 = T220 ^ 1'h1;
  assign T220 = T221 | io_in_1_valid;
  assign T221 = T222 | io_in_0_valid;
  assign T222 = T223 | T176;
  assign T223 = T224 | T179;
  assign T224 = T225 | T182;
  assign T225 = T226 | T185;
  assign T226 = T227 | T188;
  assign T227 = T228 | T191;
  assign T228 = T196 | T194;
  assign T229 = T231 & T230;
  assign T230 = last_grant < 3'h2;
  assign T231 = T232 ^ 1'h1;
  assign T232 = T196 | T194;
  assign T233 = lockIdx == 3'h2;
  assign io_in_3_ready = T234;
  assign T234 = T235 & io_out_ready;
  assign T235 = locked ? T253 : T236;
  assign T236 = T248 | T237;
  assign T237 = T238 ^ 1'h1;
  assign T238 = T239 | io_in_2_valid;
  assign T239 = T240 | io_in_1_valid;
  assign T240 = T241 | io_in_0_valid;
  assign T241 = T242 | T176;
  assign T242 = T243 | T179;
  assign T243 = T244 | T182;
  assign T244 = T245 | T185;
  assign T245 = T246 | T188;
  assign T246 = T247 | T191;
  assign T247 = T196 | T194;
  assign T248 = T250 & T249;
  assign T249 = last_grant < 3'h3;
  assign T250 = T251 ^ 1'h1;
  assign T251 = T252 | T191;
  assign T252 = T196 | T194;
  assign T253 = lockIdx == 3'h3;
  assign io_in_4_ready = T254;
  assign T254 = T255 & io_out_ready;
  assign T255 = locked ? T275 : T256;
  assign T256 = T269 | T257;
  assign T257 = T258 ^ 1'h1;
  assign T258 = T259 | io_in_3_valid;
  assign T259 = T260 | io_in_2_valid;
  assign T260 = T261 | io_in_1_valid;
  assign T261 = T262 | io_in_0_valid;
  assign T262 = T263 | T176;
  assign T263 = T264 | T179;
  assign T264 = T265 | T182;
  assign T265 = T266 | T185;
  assign T266 = T267 | T188;
  assign T267 = T268 | T191;
  assign T268 = T196 | T194;
  assign T269 = T271 & T270;
  assign T270 = last_grant < 3'h4;
  assign T271 = T272 ^ 1'h1;
  assign T272 = T273 | T188;
  assign T273 = T274 | T191;
  assign T274 = T196 | T194;
  assign T275 = lockIdx == 3'h4;
  assign io_in_5_ready = T276;
  assign T276 = T277 & io_out_ready;
  assign T277 = locked ? T299 : T278;
  assign T278 = T292 | T279;
  assign T279 = T280 ^ 1'h1;
  assign T280 = T281 | io_in_4_valid;
  assign T281 = T282 | io_in_3_valid;
  assign T282 = T283 | io_in_2_valid;
  assign T283 = T284 | io_in_1_valid;
  assign T284 = T285 | io_in_0_valid;
  assign T285 = T286 | T176;
  assign T286 = T287 | T179;
  assign T287 = T288 | T182;
  assign T288 = T289 | T185;
  assign T289 = T290 | T188;
  assign T290 = T291 | T191;
  assign T291 = T196 | T194;
  assign T292 = T294 & T293;
  assign T293 = last_grant < 3'h5;
  assign T294 = T295 ^ 1'h1;
  assign T295 = T296 | T185;
  assign T296 = T297 | T188;
  assign T297 = T298 | T191;
  assign T298 = T196 | T194;
  assign T299 = lockIdx == 3'h5;
  assign io_in_6_ready = T300;
  assign T300 = T301 & io_out_ready;
  assign T301 = locked ? T325 : T302;
  assign T302 = T317 | T303;
  assign T303 = T304 ^ 1'h1;
  assign T304 = T305 | io_in_5_valid;
  assign T305 = T306 | io_in_4_valid;
  assign T306 = T307 | io_in_3_valid;
  assign T307 = T308 | io_in_2_valid;
  assign T308 = T309 | io_in_1_valid;
  assign T309 = T310 | io_in_0_valid;
  assign T310 = T311 | T176;
  assign T311 = T312 | T179;
  assign T312 = T313 | T182;
  assign T313 = T314 | T185;
  assign T314 = T315 | T188;
  assign T315 = T316 | T191;
  assign T316 = T196 | T194;
  assign T317 = T319 & T318;
  assign T318 = last_grant < 3'h6;
  assign T319 = T320 ^ 1'h1;
  assign T320 = T321 | T182;
  assign T321 = T322 | T185;
  assign T322 = T323 | T188;
  assign T323 = T324 | T191;
  assign T324 = T196 | T194;
  assign T325 = lockIdx == 3'h6;
  assign io_in_7_ready = T326;
  assign T326 = T327 & io_out_ready;
  assign T327 = locked ? T353 : T328;
  assign T328 = T344 | T329;
  assign T329 = T330 ^ 1'h1;
  assign T330 = T331 | io_in_6_valid;
  assign T331 = T332 | io_in_5_valid;
  assign T332 = T333 | io_in_4_valid;
  assign T333 = T334 | io_in_3_valid;
  assign T334 = T335 | io_in_2_valid;
  assign T335 = T336 | io_in_1_valid;
  assign T336 = T337 | io_in_0_valid;
  assign T337 = T338 | T176;
  assign T338 = T339 | T179;
  assign T339 = T340 | T182;
  assign T340 = T341 | T185;
  assign T341 = T342 | T188;
  assign T342 = T343 | T191;
  assign T343 = T196 | T194;
  assign T344 = T346 & T345;
  assign T345 = last_grant < 3'h7;
  assign T346 = T347 ^ 1'h1;
  assign T347 = T348 | T179;
  assign T348 = T349 | T182;
  assign T349 = T350 | T185;
  assign T350 = T351 | T188;
  assign T351 = T352 | T191;
  assign T352 = T196 | T194;
  assign T353 = lockIdx == 3'h7;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T17) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h7;
    end else if(T45) begin
      lockIdx <= T31;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T53) begin
      locked <= 1'h0;
    end else if(T45) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R56 <= 2'h0;
    end else if(T47) begin
      R56 <= T55;
    end
  end
endmodule

module ClientUncachedTileLinkIOArbiter(input clk, input reset,
    output io_in_7_acquire_ready,
    input  io_in_7_acquire_valid,
    input [25:0] io_in_7_acquire_bits_addr_block,
    input [3:0] io_in_7_acquire_bits_client_xact_id,
    input [1:0] io_in_7_acquire_bits_addr_beat,
    input  io_in_7_acquire_bits_is_builtin_type,
    input [2:0] io_in_7_acquire_bits_a_type,
    input [16:0] io_in_7_acquire_bits_union,
    input [3:0] io_in_7_acquire_bits_data,
    input  io_in_7_grant_ready,
    output io_in_7_grant_valid,
    output[1:0] io_in_7_grant_bits_addr_beat,
    output[3:0] io_in_7_grant_bits_client_xact_id,
    output io_in_7_grant_bits_manager_xact_id,
    output io_in_7_grant_bits_is_builtin_type,
    output[3:0] io_in_7_grant_bits_g_type,
    output[3:0] io_in_7_grant_bits_data,
    output io_in_6_acquire_ready,
    input  io_in_6_acquire_valid,
    input [25:0] io_in_6_acquire_bits_addr_block,
    input [3:0] io_in_6_acquire_bits_client_xact_id,
    input [1:0] io_in_6_acquire_bits_addr_beat,
    input  io_in_6_acquire_bits_is_builtin_type,
    input [2:0] io_in_6_acquire_bits_a_type,
    input [16:0] io_in_6_acquire_bits_union,
    input [3:0] io_in_6_acquire_bits_data,
    input  io_in_6_grant_ready,
    output io_in_6_grant_valid,
    output[1:0] io_in_6_grant_bits_addr_beat,
    output[3:0] io_in_6_grant_bits_client_xact_id,
    output io_in_6_grant_bits_manager_xact_id,
    output io_in_6_grant_bits_is_builtin_type,
    output[3:0] io_in_6_grant_bits_g_type,
    output[3:0] io_in_6_grant_bits_data,
    output io_in_5_acquire_ready,
    input  io_in_5_acquire_valid,
    input [25:0] io_in_5_acquire_bits_addr_block,
    input [3:0] io_in_5_acquire_bits_client_xact_id,
    input [1:0] io_in_5_acquire_bits_addr_beat,
    input  io_in_5_acquire_bits_is_builtin_type,
    input [2:0] io_in_5_acquire_bits_a_type,
    input [16:0] io_in_5_acquire_bits_union,
    input [3:0] io_in_5_acquire_bits_data,
    input  io_in_5_grant_ready,
    output io_in_5_grant_valid,
    output[1:0] io_in_5_grant_bits_addr_beat,
    output[3:0] io_in_5_grant_bits_client_xact_id,
    output io_in_5_grant_bits_manager_xact_id,
    output io_in_5_grant_bits_is_builtin_type,
    output[3:0] io_in_5_grant_bits_g_type,
    output[3:0] io_in_5_grant_bits_data,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [25:0] io_in_4_acquire_bits_addr_block,
    input [3:0] io_in_4_acquire_bits_client_xact_id,
    input [1:0] io_in_4_acquire_bits_addr_beat,
    input  io_in_4_acquire_bits_is_builtin_type,
    input [2:0] io_in_4_acquire_bits_a_type,
    input [16:0] io_in_4_acquire_bits_union,
    input [3:0] io_in_4_acquire_bits_data,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_addr_beat,
    output[3:0] io_in_4_grant_bits_client_xact_id,
    output io_in_4_grant_bits_manager_xact_id,
    output io_in_4_grant_bits_is_builtin_type,
    output[3:0] io_in_4_grant_bits_g_type,
    output[3:0] io_in_4_grant_bits_data,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [25:0] io_in_3_acquire_bits_addr_block,
    input [3:0] io_in_3_acquire_bits_client_xact_id,
    input [1:0] io_in_3_acquire_bits_addr_beat,
    input  io_in_3_acquire_bits_is_builtin_type,
    input [2:0] io_in_3_acquire_bits_a_type,
    input [16:0] io_in_3_acquire_bits_union,
    input [3:0] io_in_3_acquire_bits_data,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_addr_beat,
    output[3:0] io_in_3_grant_bits_client_xact_id,
    output io_in_3_grant_bits_manager_xact_id,
    output io_in_3_grant_bits_is_builtin_type,
    output[3:0] io_in_3_grant_bits_g_type,
    output[3:0] io_in_3_grant_bits_data,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [25:0] io_in_2_acquire_bits_addr_block,
    input [3:0] io_in_2_acquire_bits_client_xact_id,
    input [1:0] io_in_2_acquire_bits_addr_beat,
    input  io_in_2_acquire_bits_is_builtin_type,
    input [2:0] io_in_2_acquire_bits_a_type,
    input [16:0] io_in_2_acquire_bits_union,
    input [3:0] io_in_2_acquire_bits_data,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_addr_beat,
    output[3:0] io_in_2_grant_bits_client_xact_id,
    output io_in_2_grant_bits_manager_xact_id,
    output io_in_2_grant_bits_is_builtin_type,
    output[3:0] io_in_2_grant_bits_g_type,
    output[3:0] io_in_2_grant_bits_data,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [25:0] io_in_1_acquire_bits_addr_block,
    input [3:0] io_in_1_acquire_bits_client_xact_id,
    input [1:0] io_in_1_acquire_bits_addr_beat,
    input  io_in_1_acquire_bits_is_builtin_type,
    input [2:0] io_in_1_acquire_bits_a_type,
    input [16:0] io_in_1_acquire_bits_union,
    input [3:0] io_in_1_acquire_bits_data,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_addr_beat,
    output[3:0] io_in_1_grant_bits_client_xact_id,
    output io_in_1_grant_bits_manager_xact_id,
    output io_in_1_grant_bits_is_builtin_type,
    output[3:0] io_in_1_grant_bits_g_type,
    output[3:0] io_in_1_grant_bits_data,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [25:0] io_in_0_acquire_bits_addr_block,
    input [3:0] io_in_0_acquire_bits_client_xact_id,
    input [1:0] io_in_0_acquire_bits_addr_beat,
    input  io_in_0_acquire_bits_is_builtin_type,
    input [2:0] io_in_0_acquire_bits_a_type,
    input [16:0] io_in_0_acquire_bits_union,
    input [3:0] io_in_0_acquire_bits_data,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_addr_beat,
    output[3:0] io_in_0_grant_bits_client_xact_id,
    output io_in_0_grant_bits_manager_xact_id,
    output io_in_0_grant_bits_is_builtin_type,
    output[3:0] io_in_0_grant_bits_g_type,
    output[3:0] io_in_0_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[3:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[3:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [3:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [3:0] io_out_grant_bits_data
);

  wire[3:0] T56;
  wire[6:0] T0;
  wire[3:0] T57;
  wire[6:0] T1;
  wire[3:0] T58;
  wire[6:0] T2;
  wire[3:0] T59;
  wire[6:0] T3;
  wire[3:0] T60;
  wire[6:0] T4;
  wire[3:0] T61;
  wire[6:0] T5;
  wire[3:0] T62;
  wire[6:0] T6;
  wire[3:0] T63;
  wire[6:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire T37;
  wire[2:0] T38;
  wire[2:0] T39;
  wire[3:0] T64;
  wire T40;
  wire T41;
  wire[3:0] T65;
  wire T42;
  wire T43;
  wire[3:0] T66;
  wire T44;
  wire T45;
  wire[3:0] T67;
  wire T46;
  wire T47;
  wire[3:0] T68;
  wire T48;
  wire T49;
  wire[3:0] T69;
  wire T50;
  wire T51;
  wire[3:0] T70;
  wire T52;
  wire T53;
  wire[3:0] T71;
  wire T54;
  wire T55;
  wire LockingRRArbiter_io_in_7_ready;
  wire LockingRRArbiter_io_in_6_ready;
  wire LockingRRArbiter_io_in_5_ready;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[25:0] LockingRRArbiter_io_out_bits_addr_block;
  wire[3:0] LockingRRArbiter_io_out_bits_client_xact_id;
  wire[1:0] LockingRRArbiter_io_out_bits_addr_beat;
  wire LockingRRArbiter_io_out_bits_is_builtin_type;
  wire[2:0] LockingRRArbiter_io_out_bits_a_type;
  wire[16:0] LockingRRArbiter_io_out_bits_union;
  wire[3:0] LockingRRArbiter_io_out_bits_data;


  assign T56 = T0[2'h3:1'h0];
  assign T0 = {io_in_0_acquire_bits_client_xact_id, 3'h0};
  assign T57 = T1[2'h3:1'h0];
  assign T1 = {io_in_1_acquire_bits_client_xact_id, 3'h1};
  assign T58 = T2[2'h3:1'h0];
  assign T2 = {io_in_2_acquire_bits_client_xact_id, 3'h2};
  assign T59 = T3[2'h3:1'h0];
  assign T3 = {io_in_3_acquire_bits_client_xact_id, 3'h3};
  assign T60 = T4[2'h3:1'h0];
  assign T4 = {io_in_4_acquire_bits_client_xact_id, 3'h4};
  assign T61 = T5[2'h3:1'h0];
  assign T5 = {io_in_5_acquire_bits_client_xact_id, 3'h5};
  assign T62 = T6[2'h3:1'h0];
  assign T6 = {io_in_6_acquire_bits_client_xact_id, 3'h6};
  assign T63 = T7[2'h3:1'h0];
  assign T7 = {io_in_7_acquire_bits_client_xact_id, 3'h7};
  assign io_out_grant_ready = T8;
  assign T8 = T37 ? io_in_7_grant_ready : T9;
  assign T9 = T34 ? io_in_6_grant_ready : T10;
  assign T10 = T31 ? io_in_5_grant_ready : T11;
  assign T11 = T28 ? io_in_4_grant_ready : T12;
  assign T12 = T25 ? io_in_3_grant_ready : T13;
  assign T13 = T22 ? io_in_2_grant_ready : T14;
  assign T14 = T19 ? io_in_1_grant_ready : T15;
  assign T15 = T16 ? io_in_0_grant_ready : 1'h0;
  assign T16 = T17 == 3'h0;
  assign T17 = T18;
  assign T18 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T19 = T20 == 3'h1;
  assign T20 = T21;
  assign T21 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T22 = T23 == 3'h2;
  assign T23 = T24;
  assign T24 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T25 = T26 == 3'h3;
  assign T26 = T27;
  assign T27 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T28 = T29 == 3'h4;
  assign T29 = T30;
  assign T30 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T31 = T32 == 3'h5;
  assign T32 = T33;
  assign T33 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T34 = T35 == 3'h6;
  assign T35 = T36;
  assign T36 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T37 = T38 == 3'h7;
  assign T38 = T39;
  assign T39 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign io_out_acquire_bits_data = LockingRRArbiter_io_out_bits_data;
  assign io_out_acquire_bits_union = LockingRRArbiter_io_out_bits_union;
  assign io_out_acquire_bits_a_type = LockingRRArbiter_io_out_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = LockingRRArbiter_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = LockingRRArbiter_io_out_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = LockingRRArbiter_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = LockingRRArbiter_io_out_bits_addr_block;
  assign io_out_acquire_valid = LockingRRArbiter_io_out_valid;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_client_xact_id = T64;
  assign T64 = {3'h0, T40};
  assign T40 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_valid = T41;
  assign T41 = T16 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = LockingRRArbiter_io_in_0_ready;
  assign io_in_1_grant_bits_data = io_out_grant_bits_data;
  assign io_in_1_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_1_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_1_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_1_grant_bits_client_xact_id = T65;
  assign T65 = {3'h0, T42};
  assign T42 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_1_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_1_grant_valid = T43;
  assign T43 = T19 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = LockingRRArbiter_io_in_1_ready;
  assign io_in_2_grant_bits_data = io_out_grant_bits_data;
  assign io_in_2_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_2_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_2_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_2_grant_bits_client_xact_id = T66;
  assign T66 = {3'h0, T44};
  assign T44 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_2_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_2_grant_valid = T45;
  assign T45 = T22 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = LockingRRArbiter_io_in_2_ready;
  assign io_in_3_grant_bits_data = io_out_grant_bits_data;
  assign io_in_3_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_3_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_3_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_3_grant_bits_client_xact_id = T67;
  assign T67 = {3'h0, T46};
  assign T46 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_3_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_3_grant_valid = T47;
  assign T47 = T25 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = LockingRRArbiter_io_in_3_ready;
  assign io_in_4_grant_bits_data = io_out_grant_bits_data;
  assign io_in_4_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_4_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_4_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_4_grant_bits_client_xact_id = T68;
  assign T68 = {3'h0, T48};
  assign T48 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_4_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_4_grant_valid = T49;
  assign T49 = T28 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = LockingRRArbiter_io_in_4_ready;
  assign io_in_5_grant_bits_data = io_out_grant_bits_data;
  assign io_in_5_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_5_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_5_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_5_grant_bits_client_xact_id = T69;
  assign T69 = {3'h0, T50};
  assign T50 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_5_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_5_grant_valid = T51;
  assign T51 = T31 ? io_out_grant_valid : 1'h0;
  assign io_in_5_acquire_ready = LockingRRArbiter_io_in_5_ready;
  assign io_in_6_grant_bits_data = io_out_grant_bits_data;
  assign io_in_6_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_6_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_6_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_6_grant_bits_client_xact_id = T70;
  assign T70 = {3'h0, T52};
  assign T52 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_6_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_6_grant_valid = T53;
  assign T53 = T34 ? io_out_grant_valid : 1'h0;
  assign io_in_6_acquire_ready = LockingRRArbiter_io_in_6_ready;
  assign io_in_7_grant_bits_data = io_out_grant_bits_data;
  assign io_in_7_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_7_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_7_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_7_grant_bits_client_xact_id = T71;
  assign T71 = {3'h0, T54};
  assign T54 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_7_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_7_grant_valid = T55;
  assign T55 = T37 ? io_out_grant_valid : 1'h0;
  assign io_in_7_acquire_ready = LockingRRArbiter_io_in_7_ready;
  LockingRRArbiter_5 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_7_ready( LockingRRArbiter_io_in_7_ready ),
       .io_in_7_valid( io_in_7_acquire_valid ),
       .io_in_7_bits_addr_block( io_in_7_acquire_bits_addr_block ),
       .io_in_7_bits_client_xact_id( T63 ),
       .io_in_7_bits_addr_beat( io_in_7_acquire_bits_addr_beat ),
       .io_in_7_bits_is_builtin_type( io_in_7_acquire_bits_is_builtin_type ),
       .io_in_7_bits_a_type( io_in_7_acquire_bits_a_type ),
       .io_in_7_bits_union( io_in_7_acquire_bits_union ),
       .io_in_7_bits_data( io_in_7_acquire_bits_data ),
       .io_in_6_ready( LockingRRArbiter_io_in_6_ready ),
       .io_in_6_valid( io_in_6_acquire_valid ),
       .io_in_6_bits_addr_block( io_in_6_acquire_bits_addr_block ),
       .io_in_6_bits_client_xact_id( T62 ),
       .io_in_6_bits_addr_beat( io_in_6_acquire_bits_addr_beat ),
       .io_in_6_bits_is_builtin_type( io_in_6_acquire_bits_is_builtin_type ),
       .io_in_6_bits_a_type( io_in_6_acquire_bits_a_type ),
       .io_in_6_bits_union( io_in_6_acquire_bits_union ),
       .io_in_6_bits_data( io_in_6_acquire_bits_data ),
       .io_in_5_ready( LockingRRArbiter_io_in_5_ready ),
       .io_in_5_valid( io_in_5_acquire_valid ),
       .io_in_5_bits_addr_block( io_in_5_acquire_bits_addr_block ),
       .io_in_5_bits_client_xact_id( T61 ),
       .io_in_5_bits_addr_beat( io_in_5_acquire_bits_addr_beat ),
       .io_in_5_bits_is_builtin_type( io_in_5_acquire_bits_is_builtin_type ),
       .io_in_5_bits_a_type( io_in_5_acquire_bits_a_type ),
       .io_in_5_bits_union( io_in_5_acquire_bits_union ),
       .io_in_5_bits_data( io_in_5_acquire_bits_data ),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_addr_block( io_in_4_acquire_bits_addr_block ),
       .io_in_4_bits_client_xact_id( T60 ),
       .io_in_4_bits_addr_beat( io_in_4_acquire_bits_addr_beat ),
       .io_in_4_bits_is_builtin_type( io_in_4_acquire_bits_is_builtin_type ),
       .io_in_4_bits_a_type( io_in_4_acquire_bits_a_type ),
       .io_in_4_bits_union( io_in_4_acquire_bits_union ),
       .io_in_4_bits_data( io_in_4_acquire_bits_data ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_addr_block( io_in_3_acquire_bits_addr_block ),
       .io_in_3_bits_client_xact_id( T59 ),
       .io_in_3_bits_addr_beat( io_in_3_acquire_bits_addr_beat ),
       .io_in_3_bits_is_builtin_type( io_in_3_acquire_bits_is_builtin_type ),
       .io_in_3_bits_a_type( io_in_3_acquire_bits_a_type ),
       .io_in_3_bits_union( io_in_3_acquire_bits_union ),
       .io_in_3_bits_data( io_in_3_acquire_bits_data ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_addr_block( io_in_2_acquire_bits_addr_block ),
       .io_in_2_bits_client_xact_id( T58 ),
       .io_in_2_bits_addr_beat( io_in_2_acquire_bits_addr_beat ),
       .io_in_2_bits_is_builtin_type( io_in_2_acquire_bits_is_builtin_type ),
       .io_in_2_bits_a_type( io_in_2_acquire_bits_a_type ),
       .io_in_2_bits_union( io_in_2_acquire_bits_union ),
       .io_in_2_bits_data( io_in_2_acquire_bits_data ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_addr_block( io_in_1_acquire_bits_addr_block ),
       .io_in_1_bits_client_xact_id( T57 ),
       .io_in_1_bits_addr_beat( io_in_1_acquire_bits_addr_beat ),
       .io_in_1_bits_is_builtin_type( io_in_1_acquire_bits_is_builtin_type ),
       .io_in_1_bits_a_type( io_in_1_acquire_bits_a_type ),
       .io_in_1_bits_union( io_in_1_acquire_bits_union ),
       .io_in_1_bits_data( io_in_1_acquire_bits_data ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_addr_block( io_in_0_acquire_bits_addr_block ),
       .io_in_0_bits_client_xact_id( T56 ),
       .io_in_0_bits_addr_beat( io_in_0_acquire_bits_addr_beat ),
       .io_in_0_bits_is_builtin_type( io_in_0_acquire_bits_is_builtin_type ),
       .io_in_0_bits_a_type( io_in_0_acquire_bits_a_type ),
       .io_in_0_bits_union( io_in_0_acquire_bits_union ),
       .io_in_0_bits_data( io_in_0_acquire_bits_data ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_addr_block( LockingRRArbiter_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( LockingRRArbiter_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( LockingRRArbiter_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( LockingRRArbiter_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( LockingRRArbiter_io_out_bits_a_type ),
       .io_out_bits_union( LockingRRArbiter_io_out_bits_union ),
       .io_out_bits_data( LockingRRArbiter_io_out_bits_data )
       //.io_chosen(  )
  );
endmodule

module L2BroadcastHub(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [127:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[127:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [127:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[127:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [127:0] io_outer_grant_bits_data
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[7:0] releaseMatches;
  wire[7:0] T6;
  wire[3:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[3:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[3:0] T293;
  wire[127:0] T294;
  wire[127:0] T295;
  wire[127:0] T296;
  wire[127:0] T297;
  wire[127:0] T298;
  wire[127:0] T299;
  wire[127:0] T300;
  wire[127:0] T301;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[1:0] T15;
  wire[1:0] T16;
  reg [1:0] rel_data_cnt;
  wire[1:0] T302;
  wire[1:0] T17;
  wire[1:0] T18;
  wire vwbdq_enq;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[2:0] T303;
  wire[2:0] T304;
  wire[2:0] T305;
  wire[2:0] T306;
  wire[2:0] T307;
  wire[2:0] T308;
  wire[2:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T28;
  wire T29;
  wire[3:0] T30;
  wire[3:0] T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T317;
  wire[1:0] T318;
  wire[1:0] T319;
  wire T320;
  wire[3:0] T34;
  reg [3:0] sdq_val;
  wire[3:0] T321;
  wire[3:0] T35;
  wire[3:0] T36;
  wire[3:0] T37;
  wire[3:0] T38;
  wire[3:0] T322;
  wire sdq_enq;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[3:0] T46;
  wire[3:0] T47;
  wire[3:0] T48;
  wire[3:0] T49;
  wire T50;
  wire[3:0] T51;
  wire[3:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T323;
  wire free_sdq;
  wire T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[3:0] T70;
  wire[1:0] T71;
  wire T72;
  wire T324;
  wire T325;
  wire T73;
  wire T74;
  wire[2:0] acquire_idx;
  wire[2:0] T326;
  wire[2:0] T327;
  wire[2:0] T328;
  wire[2:0] T329;
  wire[2:0] T330;
  wire[2:0] T331;
  wire[2:0] T332;
  wire T333;
  wire[7:0] acquireReadys;
  wire[7:0] T76;
  wire[3:0] T77;
  wire[1:0] T78;
  wire[1:0] T79;
  wire[3:0] T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire[2:0] T340;
  wire[2:0] T341;
  wire[2:0] T342;
  wire[2:0] T343;
  wire[2:0] T344;
  wire[2:0] T345;
  wire[2:0] T346;
  wire T347;
  wire[7:0] acquireMatches;
  wire[7:0] T84;
  wire[3:0] T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire[3:0] T88;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T91;
  wire T92;
  wire T93;
  wire block_acquires;
  wire T94;
  wire sdq_rdy;
  wire T95;
  wire T96;
  wire[7:0] acquireConflicts;
  wire[7:0] T97;
  wire[3:0] T98;
  wire[1:0] T99;
  wire[1:0] T100;
  wire[3:0] T101;
  wire[1:0] T102;
  wire[1:0] T103;
  wire[3:0] T104;
  wire[3:0] T105;
  wire[1:0] T106;
  wire[1:0] T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[3:0] T112;
  wire[3:0] T113;
  wire[1:0] T114;
  wire[1:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire[3:0] T120;
  wire[3:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire[3:0] T128;
  wire[3:0] T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[3:0] T136;
  wire[3:0] T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire[3:0] T144;
  wire[3:0] T145;
  wire[1:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire[3:0] T152;
  wire[3:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire[3:0] T160;
  wire[3:0] T161;
  wire[1:0] T162;
  wire[1:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire[3:0] T168;
  wire[3:0] T169;
  wire[1:0] T170;
  wire[1:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire[3:0] T176;
  wire[3:0] T177;
  wire[1:0] T178;
  wire[1:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[3:0] T184;
  wire[3:0] T185;
  wire[1:0] T186;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[1:0] T194;
  wire[1:0] T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire[3:0] T200;
  wire[3:0] T201;
  wire[1:0] T202;
  wire[1:0] T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire[3:0] T208;
  wire[3:0] T209;
  wire[1:0] T210;
  wire[1:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[127:0] T216;
  wire[127:0] T217;
  wire[127:0] T218;
  wire[127:0] T219;
  reg [127:0] vwbdq_0;
  wire[127:0] T220;
  wire T221;
  wire T222;
  wire[3:0] T223;
  wire[1:0] T224;
  reg [127:0] vwbdq_1;
  wire[127:0] T225;
  wire T226;
  wire T227;
  wire T228;
  wire[1:0] T229;
  wire[127:0] T230;
  reg [127:0] vwbdq_2;
  wire[127:0] T231;
  wire T232;
  wire T233;
  reg [127:0] vwbdq_3;
  wire[127:0] T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire[127:0] T240;
  wire[127:0] T241;
  reg [127:0] sdq_0;
  wire[127:0] T242;
  wire T243;
  wire T244;
  wire[3:0] T245;
  wire[1:0] T246;
  reg [127:0] sdq_1;
  wire[127:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[1:0] T251;
  wire[127:0] T252;
  reg [127:0] sdq_2;
  wire[127:0] T253;
  wire T254;
  wire T255;
  reg [127:0] sdq_3;
  wire[127:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire[2:0] T265;
  wire[2:0] T266;
  wire T267;
  wire[7:0] releaseReadys;
  wire[7:0] T268;
  wire[3:0] T269;
  wire[1:0] T270;
  wire[1:0] T271;
  wire[3:0] T272;
  wire[1:0] T273;
  wire[1:0] T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[2:0] T279;
  wire[2:0] T354;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready;
  wire BroadcastVoluntaryReleaseTracker_io_inner_grant_valid;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id;
  wire BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id;
  wire BroadcastVoluntaryReleaseTracker_io_inner_finish_ready;
  wire BroadcastVoluntaryReleaseTracker_io_inner_probe_valid;
  wire BroadcastVoluntaryReleaseTracker_io_inner_release_ready;
  wire BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid;
  wire[25:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat;
  wire BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data;
  wire BroadcastVoluntaryReleaseTracker_io_outer_grant_ready;
  wire BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict;
  wire BroadcastVoluntaryReleaseTracker_io_has_acquire_match;
  wire BroadcastVoluntaryReleaseTracker_io_has_release_match;
  wire BroadcastAcquireTracker_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_io_inner_finish_ready;
  wire BroadcastAcquireTracker_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_io_inner_release_ready;
  wire BroadcastAcquireTracker_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_io_outer_grant_ready;
  wire BroadcastAcquireTracker_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_io_has_acquire_match;
  wire BroadcastAcquireTracker_io_has_release_match;
  wire BroadcastAcquireTracker_1_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_1_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_1_io_inner_finish_ready;
  wire BroadcastAcquireTracker_1_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_1_io_inner_release_ready;
  wire BroadcastAcquireTracker_1_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_1_io_outer_grant_ready;
  wire BroadcastAcquireTracker_1_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_1_io_has_acquire_match;
  wire BroadcastAcquireTracker_1_io_has_release_match;
  wire BroadcastAcquireTracker_2_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_2_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_2_io_inner_finish_ready;
  wire BroadcastAcquireTracker_2_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_2_io_inner_release_ready;
  wire BroadcastAcquireTracker_2_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_2_io_outer_grant_ready;
  wire BroadcastAcquireTracker_2_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_2_io_has_acquire_match;
  wire BroadcastAcquireTracker_2_io_has_release_match;
  wire BroadcastAcquireTracker_3_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_3_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_3_io_inner_finish_ready;
  wire BroadcastAcquireTracker_3_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_3_io_inner_release_ready;
  wire BroadcastAcquireTracker_3_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_3_io_outer_grant_ready;
  wire BroadcastAcquireTracker_3_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_3_io_has_acquire_match;
  wire BroadcastAcquireTracker_3_io_has_release_match;
  wire BroadcastAcquireTracker_4_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_4_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_4_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_4_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_4_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_4_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_4_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_4_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_4_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_4_io_inner_finish_ready;
  wire BroadcastAcquireTracker_4_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_4_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_4_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_4_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_4_io_inner_release_ready;
  wire BroadcastAcquireTracker_4_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_4_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_4_io_outer_grant_ready;
  wire BroadcastAcquireTracker_4_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_4_io_has_acquire_match;
  wire BroadcastAcquireTracker_4_io_has_release_match;
  wire BroadcastAcquireTracker_5_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_5_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_5_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_5_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_5_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_5_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_5_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_5_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_5_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_5_io_inner_finish_ready;
  wire BroadcastAcquireTracker_5_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_5_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_5_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_5_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_5_io_inner_release_ready;
  wire BroadcastAcquireTracker_5_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_5_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_5_io_outer_grant_ready;
  wire BroadcastAcquireTracker_5_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_5_io_has_acquire_match;
  wire BroadcastAcquireTracker_5_io_has_release_match;
  wire BroadcastAcquireTracker_6_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_6_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_6_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_6_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_6_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_6_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_6_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_6_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_6_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_6_io_inner_finish_ready;
  wire BroadcastAcquireTracker_6_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_6_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_6_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_6_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_6_io_inner_release_ready;
  wire BroadcastAcquireTracker_6_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_6_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_6_io_outer_grant_ready;
  wire BroadcastAcquireTracker_6_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_6_io_has_acquire_match;
  wire BroadcastAcquireTracker_6_io_has_release_match;
  wire LockingRRArbiter_io_in_7_ready;
  wire LockingRRArbiter_io_in_6_ready;
  wire LockingRRArbiter_io_in_5_ready;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[1:0] LockingRRArbiter_io_out_bits_client_xact_id;
  wire[3:0] LockingRRArbiter_io_out_bits_manager_xact_id;
  wire LockingRRArbiter_io_out_bits_is_builtin_type;
  wire[3:0] LockingRRArbiter_io_out_bits_g_type;
  wire[1:0] LockingRRArbiter_io_out_bits_client_id;
  wire LockingRRArbiter_1_io_in_7_ready;
  wire LockingRRArbiter_1_io_in_6_ready;
  wire LockingRRArbiter_1_io_in_5_ready;
  wire LockingRRArbiter_1_io_in_4_ready;
  wire LockingRRArbiter_1_io_in_3_ready;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[25:0] LockingRRArbiter_1_io_out_bits_addr_block;
  wire[1:0] LockingRRArbiter_1_io_out_bits_p_type;
  wire[1:0] LockingRRArbiter_1_io_out_bits_client_id;
  wire outer_arb_io_in_7_acquire_ready;
  wire outer_arb_io_in_7_grant_valid;
  wire[1:0] outer_arb_io_in_7_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_7_grant_bits_client_xact_id;
  wire outer_arb_io_in_7_grant_bits_manager_xact_id;
  wire outer_arb_io_in_7_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_7_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_7_grant_bits_data;
  wire outer_arb_io_in_6_acquire_ready;
  wire outer_arb_io_in_6_grant_valid;
  wire[1:0] outer_arb_io_in_6_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_6_grant_bits_client_xact_id;
  wire outer_arb_io_in_6_grant_bits_manager_xact_id;
  wire outer_arb_io_in_6_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_6_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_6_grant_bits_data;
  wire outer_arb_io_in_5_acquire_ready;
  wire outer_arb_io_in_5_grant_valid;
  wire[1:0] outer_arb_io_in_5_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_5_grant_bits_client_xact_id;
  wire outer_arb_io_in_5_grant_bits_manager_xact_id;
  wire outer_arb_io_in_5_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_5_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_5_grant_bits_data;
  wire outer_arb_io_in_4_acquire_ready;
  wire outer_arb_io_in_4_grant_valid;
  wire[1:0] outer_arb_io_in_4_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_4_grant_bits_client_xact_id;
  wire outer_arb_io_in_4_grant_bits_manager_xact_id;
  wire outer_arb_io_in_4_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_4_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_4_grant_bits_data;
  wire outer_arb_io_in_3_acquire_ready;
  wire outer_arb_io_in_3_grant_valid;
  wire[1:0] outer_arb_io_in_3_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_3_grant_bits_client_xact_id;
  wire outer_arb_io_in_3_grant_bits_manager_xact_id;
  wire outer_arb_io_in_3_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_3_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_3_grant_bits_data;
  wire outer_arb_io_in_2_acquire_ready;
  wire outer_arb_io_in_2_grant_valid;
  wire[1:0] outer_arb_io_in_2_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_2_grant_bits_client_xact_id;
  wire outer_arb_io_in_2_grant_bits_manager_xact_id;
  wire outer_arb_io_in_2_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_2_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_2_grant_bits_data;
  wire outer_arb_io_in_1_acquire_ready;
  wire outer_arb_io_in_1_grant_valid;
  wire[1:0] outer_arb_io_in_1_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_1_grant_bits_client_xact_id;
  wire outer_arb_io_in_1_grant_bits_manager_xact_id;
  wire outer_arb_io_in_1_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_1_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_1_grant_bits_data;
  wire outer_arb_io_in_0_acquire_ready;
  wire outer_arb_io_in_0_grant_valid;
  wire[1:0] outer_arb_io_in_0_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_0_grant_bits_client_xact_id;
  wire outer_arb_io_in_0_grant_bits_manager_xact_id;
  wire outer_arb_io_in_0_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_0_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_0_grant_bits_data;
  wire outer_arb_io_out_acquire_valid;
  wire[25:0] outer_arb_io_out_acquire_bits_addr_block;
  wire[3:0] outer_arb_io_out_acquire_bits_client_xact_id;
  wire[1:0] outer_arb_io_out_acquire_bits_addr_beat;
  wire outer_arb_io_out_acquire_bits_is_builtin_type;
  wire[2:0] outer_arb_io_out_acquire_bits_a_type;
  wire[16:0] outer_arb_io_out_acquire_bits_union;
  wire[3:0] outer_arb_io_out_acquire_bits_data;
  wire outer_arb_io_out_grant_ready;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    rel_data_cnt = {1{$random}};
    sdq_val = {1{$random}};
    vwbdq_0 = {4{$random}};
    vwbdq_1 = {4{$random}};
    vwbdq_2 = {4{$random}};
    vwbdq_3 = {4{$random}};
    sdq_0 = {4{$random}};
    sdq_1 = {4{$random}};
    sdq_2 = {4{$random}};
    sdq_3 = {4{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_inner_release_valid & T4;
  assign T4 = T5 ^ 1'h1;
  assign T5 = releaseMatches != 8'h0;
  assign releaseMatches = T6;
  assign T6 = {T10, T7};
  assign T7 = {T9, T8};
  assign T8 = {BroadcastAcquireTracker_io_has_release_match, BroadcastVoluntaryReleaseTracker_io_has_release_match};
  assign T9 = {BroadcastAcquireTracker_2_io_has_release_match, BroadcastAcquireTracker_1_io_has_release_match};
  assign T10 = {T12, T11};
  assign T11 = {BroadcastAcquireTracker_4_io_has_release_match, BroadcastAcquireTracker_3_io_has_release_match};
  assign T12 = {BroadcastAcquireTracker_6_io_has_release_match, BroadcastAcquireTracker_5_io_has_release_match};
  assign T293 = io_outer_grant_bits_data[2'h3:1'h0];
  assign T294 = {124'h0, BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data};
  assign T295 = {124'h0, BroadcastAcquireTracker_io_inner_grant_bits_data};
  assign T296 = {124'h0, BroadcastAcquireTracker_1_io_inner_grant_bits_data};
  assign T297 = {124'h0, BroadcastAcquireTracker_2_io_inner_grant_bits_data};
  assign T298 = {124'h0, BroadcastAcquireTracker_3_io_inner_grant_bits_data};
  assign T299 = {124'h0, BroadcastAcquireTracker_4_io_inner_grant_bits_data};
  assign T300 = {124'h0, BroadcastAcquireTracker_5_io_inner_grant_bits_data};
  assign T301 = {124'h0, BroadcastAcquireTracker_6_io_inner_grant_bits_data};
  assign T13 = T14;
  assign T14 = {T16, T15};
  assign T15 = 2'h2;
  assign T16 = rel_data_cnt;
  assign T302 = reset ? 2'h0 : T17;
  assign T17 = vwbdq_enq ? T18 : rel_data_cnt;
  assign T18 = rel_data_cnt + 2'h1;
  assign vwbdq_enq = T24 & T19;
  assign T19 = T21 | T20;
  assign T20 = 3'h2 == io_inner_release_bits_r_type;
  assign T21 = T23 | T22;
  assign T22 = 3'h1 == io_inner_release_bits_r_type;
  assign T23 = 3'h0 == io_inner_release_bits_r_type;
  assign T24 = T25 & io_inner_release_bits_voluntary;
  assign T25 = io_inner_release_ready & io_inner_release_valid;
  assign T26 = io_inner_release_valid & T27;
  assign T27 = T303 == 3'h7;
  assign T303 = T316 ? 1'h0 : T304;
  assign T304 = T315 ? 1'h1 : T305;
  assign T305 = T314 ? 2'h2 : T306;
  assign T306 = T313 ? 2'h3 : T307;
  assign T307 = T312 ? 3'h4 : T308;
  assign T308 = T311 ? 3'h5 : T309;
  assign T309 = T310 ? 3'h6 : 3'h7;
  assign T310 = releaseMatches[3'h6:3'h6];
  assign T311 = releaseMatches[3'h5:3'h5];
  assign T312 = releaseMatches[3'h4:3'h4];
  assign T313 = releaseMatches[2'h3:2'h3];
  assign T314 = releaseMatches[2'h2:2'h2];
  assign T315 = releaseMatches[1'h1:1'h1];
  assign T316 = releaseMatches[1'h0:1'h0];
  assign T28 = io_inner_finish_valid & T29;
  assign T29 = io_inner_finish_bits_manager_xact_id == 4'h7;
  assign T30 = T31;
  assign T31 = {T33, T32};
  assign T32 = 2'h0;
  assign T33 = T317;
  assign T317 = T325 ? 1'h0 : T318;
  assign T318 = T324 ? 1'h1 : T319;
  assign T319 = T320 ? 2'h2 : 2'h3;
  assign T320 = T34[2'h2:2'h2];
  assign T34 = ~ sdq_val;
  assign T321 = reset ? 4'h0 : T35;
  assign T35 = T72 ? T36 : sdq_val;
  assign T36 = T56 | T37;
  assign T37 = T46 & T38;
  assign T38 = 4'h0 - T322;
  assign T322 = {3'h0, sdq_enq};
  assign sdq_enq = T45 & T39;
  assign T39 = io_inner_acquire_bits_is_builtin_type & T40;
  assign T40 = T42 | T41;
  assign T41 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T42 = T44 | T43;
  assign T43 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T44 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T45 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T46 = T55 ? 4'h1 : T47;
  assign T47 = T54 ? 4'h2 : T48;
  assign T48 = T53 ? 4'h4 : T49;
  assign T49 = T50 ? 4'h8 : 4'h0;
  assign T50 = T51[2'h3:2'h3];
  assign T51 = ~ T52;
  assign T52 = sdq_val[2'h3:1'h0];
  assign T53 = T51[2'h2:2'h2];
  assign T54 = T51[1'h1:1'h1];
  assign T55 = T51[1'h0:1'h0];
  assign T56 = sdq_val & T57;
  assign T57 = ~ T58;
  assign T58 = T70 & T59;
  assign T59 = 4'h0 - T323;
  assign T323 = {3'h0, free_sdq};
  assign free_sdq = T62 & T60;
  assign T60 = T61 == 2'h0;
  assign T61 = outer_arb_io_out_acquire_bits_data[1'h1:1'h0];
  assign T62 = T69 & T63;
  assign T63 = io_outer_acquire_bits_is_builtin_type & T64;
  assign T64 = T66 | T65;
  assign T65 = 3'h4 == io_outer_acquire_bits_a_type;
  assign T66 = T68 | T67;
  assign T67 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T68 = 3'h2 == io_outer_acquire_bits_a_type;
  assign T69 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T70 = 1'h1 << T71;
  assign T71 = outer_arb_io_out_acquire_bits_data[2'h3:2'h2];
  assign T72 = io_outer_acquire_valid | sdq_enq;
  assign T324 = T34[1'h1:1'h1];
  assign T325 = T34[1'h0:1'h0];
  assign T73 = T92 & T74;
  assign T74 = acquire_idx == 3'h7;
  assign acquire_idx = T91 ? T340 : T326;
  assign T326 = T339 ? 1'h0 : T327;
  assign T327 = T338 ? 1'h1 : T328;
  assign T328 = T337 ? 2'h2 : T329;
  assign T329 = T336 ? 2'h3 : T330;
  assign T330 = T335 ? 3'h4 : T331;
  assign T331 = T334 ? 3'h5 : T332;
  assign T332 = T333 ? 3'h6 : 3'h7;
  assign T333 = acquireReadys[3'h6:3'h6];
  assign acquireReadys = T76;
  assign T76 = {T80, T77};
  assign T77 = {T79, T78};
  assign T78 = {BroadcastAcquireTracker_io_inner_acquire_ready, BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready};
  assign T79 = {BroadcastAcquireTracker_2_io_inner_acquire_ready, BroadcastAcquireTracker_1_io_inner_acquire_ready};
  assign T80 = {T82, T81};
  assign T81 = {BroadcastAcquireTracker_4_io_inner_acquire_ready, BroadcastAcquireTracker_3_io_inner_acquire_ready};
  assign T82 = {BroadcastAcquireTracker_6_io_inner_acquire_ready, BroadcastAcquireTracker_5_io_inner_acquire_ready};
  assign T334 = acquireReadys[3'h5:3'h5];
  assign T335 = acquireReadys[3'h4:3'h4];
  assign T336 = acquireReadys[2'h3:2'h3];
  assign T337 = acquireReadys[2'h2:2'h2];
  assign T338 = acquireReadys[1'h1:1'h1];
  assign T339 = acquireReadys[1'h0:1'h0];
  assign T340 = T353 ? 1'h0 : T341;
  assign T341 = T352 ? 1'h1 : T342;
  assign T342 = T351 ? 2'h2 : T343;
  assign T343 = T350 ? 2'h3 : T344;
  assign T344 = T349 ? 3'h4 : T345;
  assign T345 = T348 ? 3'h5 : T346;
  assign T346 = T347 ? 3'h6 : 3'h7;
  assign T347 = acquireMatches[3'h6:3'h6];
  assign acquireMatches = T84;
  assign T84 = {T88, T85};
  assign T85 = {T87, T86};
  assign T86 = {BroadcastAcquireTracker_io_has_acquire_match, BroadcastVoluntaryReleaseTracker_io_has_acquire_match};
  assign T87 = {BroadcastAcquireTracker_2_io_has_acquire_match, BroadcastAcquireTracker_1_io_has_acquire_match};
  assign T88 = {T90, T89};
  assign T89 = {BroadcastAcquireTracker_4_io_has_acquire_match, BroadcastAcquireTracker_3_io_has_acquire_match};
  assign T90 = {BroadcastAcquireTracker_6_io_has_acquire_match, BroadcastAcquireTracker_5_io_has_acquire_match};
  assign T348 = acquireMatches[3'h5:3'h5];
  assign T349 = acquireMatches[3'h4:3'h4];
  assign T350 = acquireMatches[2'h3:2'h3];
  assign T351 = acquireMatches[2'h2:2'h2];
  assign T352 = acquireMatches[1'h1:1'h1];
  assign T353 = acquireMatches[1'h0:1'h0];
  assign T91 = acquireMatches != 8'h0;
  assign T92 = io_inner_acquire_valid & T93;
  assign T93 = block_acquires ^ 1'h1;
  assign block_acquires = T96 | T94;
  assign T94 = sdq_rdy ^ 1'h1;
  assign sdq_rdy = T95 ^ 1'h1;
  assign T95 = sdq_val == 4'hf;
  assign T96 = acquireConflicts != 8'h0;
  assign acquireConflicts = T97;
  assign T97 = {T101, T98};
  assign T98 = {T100, T99};
  assign T99 = {BroadcastAcquireTracker_io_has_acquire_conflict, BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict};
  assign T100 = {BroadcastAcquireTracker_2_io_has_acquire_conflict, BroadcastAcquireTracker_1_io_has_acquire_conflict};
  assign T101 = {T103, T102};
  assign T102 = {BroadcastAcquireTracker_4_io_has_acquire_conflict, BroadcastAcquireTracker_3_io_has_acquire_conflict};
  assign T103 = {BroadcastAcquireTracker_6_io_has_acquire_conflict, BroadcastAcquireTracker_5_io_has_acquire_conflict};
  assign T104 = T105;
  assign T105 = {T107, T106};
  assign T106 = 2'h2;
  assign T107 = rel_data_cnt;
  assign T108 = io_inner_release_valid & T109;
  assign T109 = T303 == 3'h6;
  assign T110 = io_inner_finish_valid & T111;
  assign T111 = io_inner_finish_bits_manager_xact_id == 4'h6;
  assign T112 = T113;
  assign T113 = {T115, T114};
  assign T114 = 2'h0;
  assign T115 = T317;
  assign T116 = T118 & T117;
  assign T117 = acquire_idx == 3'h6;
  assign T118 = io_inner_acquire_valid & T119;
  assign T119 = block_acquires ^ 1'h1;
  assign T120 = T121;
  assign T121 = {T123, T122};
  assign T122 = 2'h2;
  assign T123 = rel_data_cnt;
  assign T124 = io_inner_release_valid & T125;
  assign T125 = T303 == 3'h5;
  assign T126 = io_inner_finish_valid & T127;
  assign T127 = io_inner_finish_bits_manager_xact_id == 4'h5;
  assign T128 = T129;
  assign T129 = {T131, T130};
  assign T130 = 2'h0;
  assign T131 = T317;
  assign T132 = T134 & T133;
  assign T133 = acquire_idx == 3'h5;
  assign T134 = io_inner_acquire_valid & T135;
  assign T135 = block_acquires ^ 1'h1;
  assign T136 = T137;
  assign T137 = {T139, T138};
  assign T138 = 2'h2;
  assign T139 = rel_data_cnt;
  assign T140 = io_inner_release_valid & T141;
  assign T141 = T303 == 3'h4;
  assign T142 = io_inner_finish_valid & T143;
  assign T143 = io_inner_finish_bits_manager_xact_id == 4'h4;
  assign T144 = T145;
  assign T145 = {T147, T146};
  assign T146 = 2'h0;
  assign T147 = T317;
  assign T148 = T150 & T149;
  assign T149 = acquire_idx == 3'h4;
  assign T150 = io_inner_acquire_valid & T151;
  assign T151 = block_acquires ^ 1'h1;
  assign T152 = T153;
  assign T153 = {T155, T154};
  assign T154 = 2'h2;
  assign T155 = rel_data_cnt;
  assign T156 = io_inner_release_valid & T157;
  assign T157 = T303 == 3'h3;
  assign T158 = io_inner_finish_valid & T159;
  assign T159 = io_inner_finish_bits_manager_xact_id == 4'h3;
  assign T160 = T161;
  assign T161 = {T163, T162};
  assign T162 = 2'h0;
  assign T163 = T317;
  assign T164 = T166 & T165;
  assign T165 = acquire_idx == 3'h3;
  assign T166 = io_inner_acquire_valid & T167;
  assign T167 = block_acquires ^ 1'h1;
  assign T168 = T169;
  assign T169 = {T171, T170};
  assign T170 = 2'h2;
  assign T171 = rel_data_cnt;
  assign T172 = io_inner_release_valid & T173;
  assign T173 = T303 == 3'h2;
  assign T174 = io_inner_finish_valid & T175;
  assign T175 = io_inner_finish_bits_manager_xact_id == 4'h2;
  assign T176 = T177;
  assign T177 = {T179, T178};
  assign T178 = 2'h0;
  assign T179 = T317;
  assign T180 = T182 & T181;
  assign T181 = acquire_idx == 3'h2;
  assign T182 = io_inner_acquire_valid & T183;
  assign T183 = block_acquires ^ 1'h1;
  assign T184 = T185;
  assign T185 = {T187, T186};
  assign T186 = 2'h2;
  assign T187 = rel_data_cnt;
  assign T188 = io_inner_release_valid & T189;
  assign T189 = T303 == 3'h1;
  assign T190 = io_inner_finish_valid & T191;
  assign T191 = io_inner_finish_bits_manager_xact_id == 4'h1;
  assign T192 = T193;
  assign T193 = {T195, T194};
  assign T194 = 2'h0;
  assign T195 = T317;
  assign T196 = T198 & T197;
  assign T197 = acquire_idx == 3'h1;
  assign T198 = io_inner_acquire_valid & T199;
  assign T199 = block_acquires ^ 1'h1;
  assign T200 = T201;
  assign T201 = {T203, T202};
  assign T202 = 2'h1;
  assign T203 = rel_data_cnt;
  assign T204 = io_inner_release_valid & T205;
  assign T205 = T303 == 3'h0;
  assign T206 = io_inner_finish_valid & T207;
  assign T207 = io_inner_finish_bits_manager_xact_id == 4'h0;
  assign T208 = T209;
  assign T209 = {T211, T210};
  assign T210 = 2'h0;
  assign T211 = T317;
  assign T212 = T214 & T213;
  assign T213 = acquire_idx == 3'h0;
  assign T214 = io_inner_acquire_valid & T215;
  assign T215 = block_acquires ^ 1'h1;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_data = T216;
  assign T216 = T261 ? T240 : T217;
  assign T217 = T239 ? T218 : io_inner_release_bits_data;
  assign T218 = T238 ? T230 : T219;
  assign T219 = T228 ? vwbdq_1 : vwbdq_0;
  assign T220 = T221 ? io_inner_release_bits_data : vwbdq_0;
  assign T221 = vwbdq_enq & T222;
  assign T222 = T223[1'h0:1'h0];
  assign T223 = 1'h1 << T224;
  assign T224 = rel_data_cnt;
  assign T225 = T226 ? io_inner_release_bits_data : vwbdq_1;
  assign T226 = vwbdq_enq & T227;
  assign T227 = T223[1'h1:1'h1];
  assign T228 = T229[1'h0:1'h0];
  assign T229 = T71;
  assign T230 = T237 ? vwbdq_3 : vwbdq_2;
  assign T231 = T232 ? io_inner_release_bits_data : vwbdq_2;
  assign T232 = vwbdq_enq & T233;
  assign T233 = T223[2'h2:2'h2];
  assign T234 = T235 ? io_inner_release_bits_data : vwbdq_3;
  assign T235 = vwbdq_enq & T236;
  assign T236 = T223[2'h3:2'h3];
  assign T237 = T229[1'h0:1'h0];
  assign T238 = T229[1'h1:1'h1];
  assign T239 = T61 == 2'h1;
  assign T240 = T260 ? T252 : T241;
  assign T241 = T250 ? sdq_1 : sdq_0;
  assign T242 = T243 ? io_inner_acquire_bits_data : sdq_0;
  assign T243 = sdq_enq & T244;
  assign T244 = T245[1'h0:1'h0];
  assign T245 = 1'h1 << T246;
  assign T246 = T317;
  assign T247 = T248 ? io_inner_acquire_bits_data : sdq_1;
  assign T248 = sdq_enq & T249;
  assign T249 = T245[1'h1:1'h1];
  assign T250 = T251[1'h0:1'h0];
  assign T251 = T71;
  assign T252 = T259 ? sdq_3 : sdq_2;
  assign T253 = T254 ? io_inner_acquire_bits_data : sdq_2;
  assign T254 = sdq_enq & T255;
  assign T255 = T245[2'h2:2'h2];
  assign T256 = T257 ? io_inner_acquire_bits_data : sdq_3;
  assign T257 = sdq_enq & T258;
  assign T258 = T245[2'h3:2'h3];
  assign T259 = T251[1'h0:1'h0];
  assign T260 = T251[1'h1:1'h1];
  assign T261 = T61 == 2'h0;
  assign io_outer_acquire_bits_union = outer_arb_io_out_acquire_bits_union;
  assign io_outer_acquire_bits_a_type = outer_arb_io_out_acquire_bits_a_type;
  assign io_outer_acquire_bits_is_builtin_type = outer_arb_io_out_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_addr_beat = outer_arb_io_out_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = outer_arb_io_out_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_block = outer_arb_io_out_acquire_bits_addr_block;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T262;
  assign T262 = T267 & T263;
  assign T263 = T264 - 1'h1;
  assign T264 = 1'h1 << T265;
  assign T265 = T266 + 3'h1;
  assign T266 = T303 - T303;
  assign T267 = releaseReadys >> T303;
  assign releaseReadys = T268;
  assign T268 = {T272, T269};
  assign T269 = {T271, T270};
  assign T270 = {BroadcastAcquireTracker_io_inner_release_ready, BroadcastVoluntaryReleaseTracker_io_inner_release_ready};
  assign T271 = {BroadcastAcquireTracker_2_io_inner_release_ready, BroadcastAcquireTracker_1_io_inner_release_ready};
  assign T272 = {T274, T273};
  assign T273 = {BroadcastAcquireTracker_4_io_inner_release_ready, BroadcastAcquireTracker_3_io_inner_release_ready};
  assign T274 = {BroadcastAcquireTracker_6_io_inner_release_ready, BroadcastAcquireTracker_5_io_inner_release_ready};
  assign io_inner_probe_bits_client_id = LockingRRArbiter_1_io_out_bits_client_id;
  assign io_inner_probe_bits_p_type = LockingRRArbiter_1_io_out_bits_p_type;
  assign io_inner_probe_bits_addr_block = LockingRRArbiter_1_io_out_bits_addr_block;
  assign io_inner_probe_valid = LockingRRArbiter_1_io_out_valid;
  assign io_inner_finish_ready = T275;
  assign T275 = T289 ? T283 : T276;
  assign T276 = T282 ? T280 : T277;
  assign T277 = T278 ? BroadcastAcquireTracker_io_inner_finish_ready : BroadcastVoluntaryReleaseTracker_io_inner_finish_ready;
  assign T278 = T279[1'h0:1'h0];
  assign T279 = T354;
  assign T354 = io_inner_finish_bits_manager_xact_id[2'h2:1'h0];
  assign T280 = T281 ? BroadcastAcquireTracker_2_io_inner_finish_ready : BroadcastAcquireTracker_1_io_inner_finish_ready;
  assign T281 = T279[1'h0:1'h0];
  assign T282 = T279[1'h1:1'h1];
  assign T283 = T288 ? T286 : T284;
  assign T284 = T285 ? BroadcastAcquireTracker_4_io_inner_finish_ready : BroadcastAcquireTracker_3_io_inner_finish_ready;
  assign T285 = T279[1'h0:1'h0];
  assign T286 = T287 ? BroadcastAcquireTracker_6_io_inner_finish_ready : BroadcastAcquireTracker_5_io_inner_finish_ready;
  assign T287 = T279[1'h0:1'h0];
  assign T288 = T279[1'h1:1'h1];
  assign T289 = T279[2'h2:2'h2];
  assign io_inner_grant_bits_client_id = LockingRRArbiter_io_out_bits_client_id;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_g_type = LockingRRArbiter_io_out_bits_g_type;
  assign io_inner_grant_bits_is_builtin_type = LockingRRArbiter_io_out_bits_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = LockingRRArbiter_io_out_bits_manager_xact_id;
  assign io_inner_grant_bits_client_xact_id = LockingRRArbiter_io_out_bits_client_xact_id;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_valid = LockingRRArbiter_io_out_valid;
  assign io_inner_acquire_ready = T290;
  assign T290 = T292 & T291;
  assign T291 = block_acquires ^ 1'h1;
  assign T292 = acquireReadys != 8'h0;
  BroadcastVoluntaryReleaseTracker BroadcastVoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T212 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T208 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_0_ready ),
       .io_inner_grant_valid( BroadcastVoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastVoluntaryReleaseTracker_io_inner_finish_ready ),
       .io_inner_finish_valid( T206 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_inner_probe_valid( BroadcastVoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_addr_block(  )
       //.io_inner_probe_bits_p_type(  )
       //.io_inner_probe_bits_client_id(  )
       .io_inner_release_ready( BroadcastVoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( T204 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_data( T200 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastVoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_0_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_0_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_0_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_0_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_0_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_0_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastVoluntaryReleaseTracker_io_has_acquire_match ),
       .io_has_release_match( BroadcastVoluntaryReleaseTracker_io_has_release_match )
  );
  BroadcastAcquireTracker_0 BroadcastAcquireTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T196 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T192 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_1_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_io_inner_finish_ready ),
       .io_inner_finish_valid( T190 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_io_inner_release_ready ),
       .io_inner_release_valid( T188 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_data( T184 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_1_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_1_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_1_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_1_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_1_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_1_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_io_has_release_match )
  );
  BroadcastAcquireTracker_1 BroadcastAcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T180 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T176 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_2_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_1_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_1_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_1_io_inner_finish_ready ),
       .io_inner_finish_valid( T174 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_1_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_1_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( T172 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_data( T168 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_1_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_1_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_1_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_2_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_2_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_2_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_2_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_2_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_2_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_1_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_1_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_1_io_has_release_match )
  );
  BroadcastAcquireTracker_2 BroadcastAcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T164 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T160 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_3_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_2_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_2_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_2_io_inner_finish_ready ),
       .io_inner_finish_valid( T158 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_2_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_2_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( T156 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_data( T152 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_2_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_2_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_2_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_3_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_3_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_3_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_3_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_3_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_3_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_2_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_2_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_2_io_has_release_match )
  );
  BroadcastAcquireTracker_3 BroadcastAcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T148 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T144 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_4_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_3_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_3_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_3_io_inner_finish_ready ),
       .io_inner_finish_valid( T142 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_3_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_3_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( T140 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_data( T136 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_3_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_3_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_3_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_4_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_4_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_4_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_4_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_4_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_4_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_3_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_3_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_3_io_has_release_match )
  );
  BroadcastAcquireTracker_4 BroadcastAcquireTracker_4(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_4_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T132 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T128 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_5_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_4_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_4_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_4_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_4_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_4_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_4_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_4_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_4_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_4_io_inner_finish_ready ),
       .io_inner_finish_valid( T126 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_5_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_4_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_4_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_4_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_4_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_4_io_inner_release_ready ),
       .io_inner_release_valid( T124 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_data( T120 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_4_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_4_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_4_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_4_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_4_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_4_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_4_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_5_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_5_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_5_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_5_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_5_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_5_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_4_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_4_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_4_io_has_release_match )
  );
  BroadcastAcquireTracker_5 BroadcastAcquireTracker_5(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_5_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T116 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T112 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_6_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_5_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_5_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_5_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_5_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_5_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_5_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_5_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_5_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_5_io_inner_finish_ready ),
       .io_inner_finish_valid( T110 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_6_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_5_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_5_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_5_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_5_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_5_io_inner_release_ready ),
       .io_inner_release_valid( T108 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_data( T104 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_5_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_5_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_5_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_5_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_5_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_5_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_5_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_6_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_6_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_6_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_6_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_6_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_6_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_5_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_5_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_5_io_has_release_match )
  );
  BroadcastAcquireTracker_6 BroadcastAcquireTracker_6(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_6_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T73 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T30 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_7_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_6_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_6_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_6_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_6_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_6_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_6_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_6_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_6_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_6_io_inner_finish_ready ),
       .io_inner_finish_valid( T28 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_7_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_6_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_6_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_6_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_6_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_6_io_inner_release_ready ),
       .io_inner_release_valid( T26 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_data( T13 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_6_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_6_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_6_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_6_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_6_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_6_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_6_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_7_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_7_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_7_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_7_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_7_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_7_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_6_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_6_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_6_io_has_release_match )
  );
  LockingRRArbiter_2 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_7_ready( LockingRRArbiter_io_in_7_ready ),
       .io_in_7_valid( BroadcastAcquireTracker_6_io_inner_grant_valid ),
       .io_in_7_bits_addr_beat( BroadcastAcquireTracker_6_io_inner_grant_bits_addr_beat ),
       .io_in_7_bits_client_xact_id( BroadcastAcquireTracker_6_io_inner_grant_bits_client_xact_id ),
       .io_in_7_bits_manager_xact_id( BroadcastAcquireTracker_6_io_inner_grant_bits_manager_xact_id ),
       .io_in_7_bits_is_builtin_type( BroadcastAcquireTracker_6_io_inner_grant_bits_is_builtin_type ),
       .io_in_7_bits_g_type( BroadcastAcquireTracker_6_io_inner_grant_bits_g_type ),
       .io_in_7_bits_data( T301 ),
       .io_in_7_bits_client_id( BroadcastAcquireTracker_6_io_inner_grant_bits_client_id ),
       .io_in_6_ready( LockingRRArbiter_io_in_6_ready ),
       .io_in_6_valid( BroadcastAcquireTracker_5_io_inner_grant_valid ),
       .io_in_6_bits_addr_beat( BroadcastAcquireTracker_5_io_inner_grant_bits_addr_beat ),
       .io_in_6_bits_client_xact_id( BroadcastAcquireTracker_5_io_inner_grant_bits_client_xact_id ),
       .io_in_6_bits_manager_xact_id( BroadcastAcquireTracker_5_io_inner_grant_bits_manager_xact_id ),
       .io_in_6_bits_is_builtin_type( BroadcastAcquireTracker_5_io_inner_grant_bits_is_builtin_type ),
       .io_in_6_bits_g_type( BroadcastAcquireTracker_5_io_inner_grant_bits_g_type ),
       .io_in_6_bits_data( T300 ),
       .io_in_6_bits_client_id( BroadcastAcquireTracker_5_io_inner_grant_bits_client_id ),
       .io_in_5_ready( LockingRRArbiter_io_in_5_ready ),
       .io_in_5_valid( BroadcastAcquireTracker_4_io_inner_grant_valid ),
       .io_in_5_bits_addr_beat( BroadcastAcquireTracker_4_io_inner_grant_bits_addr_beat ),
       .io_in_5_bits_client_xact_id( BroadcastAcquireTracker_4_io_inner_grant_bits_client_xact_id ),
       .io_in_5_bits_manager_xact_id( BroadcastAcquireTracker_4_io_inner_grant_bits_manager_xact_id ),
       .io_in_5_bits_is_builtin_type( BroadcastAcquireTracker_4_io_inner_grant_bits_is_builtin_type ),
       .io_in_5_bits_g_type( BroadcastAcquireTracker_4_io_inner_grant_bits_g_type ),
       .io_in_5_bits_data( T299 ),
       .io_in_5_bits_client_id( BroadcastAcquireTracker_4_io_inner_grant_bits_client_id ),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( BroadcastAcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_addr_beat( BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat ),
       .io_in_4_bits_client_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id ),
       .io_in_4_bits_manager_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id ),
       .io_in_4_bits_is_builtin_type( BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type ),
       .io_in_4_bits_g_type( BroadcastAcquireTracker_3_io_inner_grant_bits_g_type ),
       .io_in_4_bits_data( T298 ),
       .io_in_4_bits_client_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_id ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( BroadcastAcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_addr_beat( BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat ),
       .io_in_3_bits_client_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id ),
       .io_in_3_bits_manager_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id ),
       .io_in_3_bits_is_builtin_type( BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type ),
       .io_in_3_bits_g_type( BroadcastAcquireTracker_2_io_inner_grant_bits_g_type ),
       .io_in_3_bits_data( T297 ),
       .io_in_3_bits_client_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_id ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( BroadcastAcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_addr_beat( BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat ),
       .io_in_2_bits_client_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id ),
       .io_in_2_bits_manager_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id ),
       .io_in_2_bits_is_builtin_type( BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type ),
       .io_in_2_bits_g_type( BroadcastAcquireTracker_1_io_inner_grant_bits_g_type ),
       .io_in_2_bits_data( T296 ),
       .io_in_2_bits_client_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_id ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( BroadcastAcquireTracker_io_inner_grant_valid ),
       .io_in_1_bits_addr_beat( BroadcastAcquireTracker_io_inner_grant_bits_addr_beat ),
       .io_in_1_bits_client_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id ),
       .io_in_1_bits_manager_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id ),
       .io_in_1_bits_is_builtin_type( BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type ),
       .io_in_1_bits_g_type( BroadcastAcquireTracker_io_inner_grant_bits_g_type ),
       .io_in_1_bits_data( T295 ),
       .io_in_1_bits_client_id( BroadcastAcquireTracker_io_inner_grant_bits_client_id ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( BroadcastVoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat ),
       .io_in_0_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id ),
       .io_in_0_bits_manager_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id ),
       .io_in_0_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type ),
       .io_in_0_bits_g_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type ),
       .io_in_0_bits_data( T294 ),
       .io_in_0_bits_client_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       //.io_out_bits_addr_beat(  )
       .io_out_bits_client_xact_id( LockingRRArbiter_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( LockingRRArbiter_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( LockingRRArbiter_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( LockingRRArbiter_io_out_bits_g_type ),
       //.io_out_bits_data(  )
       .io_out_bits_client_id( LockingRRArbiter_io_out_bits_client_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_7_ready( LockingRRArbiter_1_io_in_7_ready ),
       .io_in_7_valid( BroadcastAcquireTracker_6_io_inner_probe_valid ),
       .io_in_7_bits_addr_block( BroadcastAcquireTracker_6_io_inner_probe_bits_addr_block ),
       .io_in_7_bits_p_type( BroadcastAcquireTracker_6_io_inner_probe_bits_p_type ),
       .io_in_7_bits_client_id( BroadcastAcquireTracker_6_io_inner_probe_bits_client_id ),
       .io_in_6_ready( LockingRRArbiter_1_io_in_6_ready ),
       .io_in_6_valid( BroadcastAcquireTracker_5_io_inner_probe_valid ),
       .io_in_6_bits_addr_block( BroadcastAcquireTracker_5_io_inner_probe_bits_addr_block ),
       .io_in_6_bits_p_type( BroadcastAcquireTracker_5_io_inner_probe_bits_p_type ),
       .io_in_6_bits_client_id( BroadcastAcquireTracker_5_io_inner_probe_bits_client_id ),
       .io_in_5_ready( LockingRRArbiter_1_io_in_5_ready ),
       .io_in_5_valid( BroadcastAcquireTracker_4_io_inner_probe_valid ),
       .io_in_5_bits_addr_block( BroadcastAcquireTracker_4_io_inner_probe_bits_addr_block ),
       .io_in_5_bits_p_type( BroadcastAcquireTracker_4_io_inner_probe_bits_p_type ),
       .io_in_5_bits_client_id( BroadcastAcquireTracker_4_io_inner_probe_bits_client_id ),
       .io_in_4_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( BroadcastAcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_addr_block( BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block ),
       .io_in_4_bits_p_type( BroadcastAcquireTracker_3_io_inner_probe_bits_p_type ),
       .io_in_4_bits_client_id( BroadcastAcquireTracker_3_io_inner_probe_bits_client_id ),
       .io_in_3_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( BroadcastAcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_addr_block( BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block ),
       .io_in_3_bits_p_type( BroadcastAcquireTracker_2_io_inner_probe_bits_p_type ),
       .io_in_3_bits_client_id( BroadcastAcquireTracker_2_io_inner_probe_bits_client_id ),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( BroadcastAcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_addr_block( BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block ),
       .io_in_2_bits_p_type( BroadcastAcquireTracker_1_io_inner_probe_bits_p_type ),
       .io_in_2_bits_client_id( BroadcastAcquireTracker_1_io_inner_probe_bits_client_id ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( BroadcastAcquireTracker_io_inner_probe_valid ),
       .io_in_1_bits_addr_block( BroadcastAcquireTracker_io_inner_probe_bits_addr_block ),
       .io_in_1_bits_p_type( BroadcastAcquireTracker_io_inner_probe_bits_p_type ),
       .io_in_1_bits_client_id( BroadcastAcquireTracker_io_inner_probe_bits_client_id ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( BroadcastVoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_addr_block(  )
       //.io_in_0_bits_p_type(  )
       //.io_in_0_bits_client_id(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_addr_block( LockingRRArbiter_1_io_out_bits_addr_block ),
       .io_out_bits_p_type( LockingRRArbiter_1_io_out_bits_p_type ),
       .io_out_bits_client_id( LockingRRArbiter_1_io_out_bits_client_id )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign LockingRRArbiter_1.io_in_0_bits_addr_block = {1{$random}};
    assign LockingRRArbiter_1.io_in_0_bits_p_type = {1{$random}};
    assign LockingRRArbiter_1.io_in_0_bits_client_id = {1{$random}};
// synthesis translate_on
`endif
  ClientUncachedTileLinkIOArbiter outer_arb(.clk(clk), .reset(reset),
       .io_in_7_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_in_7_acquire_valid( BroadcastAcquireTracker_6_io_outer_acquire_valid ),
       .io_in_7_acquire_bits_addr_block( BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_block ),
       .io_in_7_acquire_bits_client_xact_id( BroadcastAcquireTracker_6_io_outer_acquire_bits_client_xact_id ),
       .io_in_7_acquire_bits_addr_beat( BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_beat ),
       .io_in_7_acquire_bits_is_builtin_type( BroadcastAcquireTracker_6_io_outer_acquire_bits_is_builtin_type ),
       .io_in_7_acquire_bits_a_type( BroadcastAcquireTracker_6_io_outer_acquire_bits_a_type ),
       .io_in_7_acquire_bits_union( BroadcastAcquireTracker_6_io_outer_acquire_bits_union ),
       .io_in_7_acquire_bits_data( BroadcastAcquireTracker_6_io_outer_acquire_bits_data ),
       .io_in_7_grant_ready( BroadcastAcquireTracker_6_io_outer_grant_ready ),
       .io_in_7_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_in_7_grant_bits_addr_beat( outer_arb_io_in_7_grant_bits_addr_beat ),
       .io_in_7_grant_bits_client_xact_id( outer_arb_io_in_7_grant_bits_client_xact_id ),
       .io_in_7_grant_bits_manager_xact_id( outer_arb_io_in_7_grant_bits_manager_xact_id ),
       .io_in_7_grant_bits_is_builtin_type( outer_arb_io_in_7_grant_bits_is_builtin_type ),
       .io_in_7_grant_bits_g_type( outer_arb_io_in_7_grant_bits_g_type ),
       .io_in_7_grant_bits_data( outer_arb_io_in_7_grant_bits_data ),
       .io_in_6_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_in_6_acquire_valid( BroadcastAcquireTracker_5_io_outer_acquire_valid ),
       .io_in_6_acquire_bits_addr_block( BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_block ),
       .io_in_6_acquire_bits_client_xact_id( BroadcastAcquireTracker_5_io_outer_acquire_bits_client_xact_id ),
       .io_in_6_acquire_bits_addr_beat( BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_beat ),
       .io_in_6_acquire_bits_is_builtin_type( BroadcastAcquireTracker_5_io_outer_acquire_bits_is_builtin_type ),
       .io_in_6_acquire_bits_a_type( BroadcastAcquireTracker_5_io_outer_acquire_bits_a_type ),
       .io_in_6_acquire_bits_union( BroadcastAcquireTracker_5_io_outer_acquire_bits_union ),
       .io_in_6_acquire_bits_data( BroadcastAcquireTracker_5_io_outer_acquire_bits_data ),
       .io_in_6_grant_ready( BroadcastAcquireTracker_5_io_outer_grant_ready ),
       .io_in_6_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_in_6_grant_bits_addr_beat( outer_arb_io_in_6_grant_bits_addr_beat ),
       .io_in_6_grant_bits_client_xact_id( outer_arb_io_in_6_grant_bits_client_xact_id ),
       .io_in_6_grant_bits_manager_xact_id( outer_arb_io_in_6_grant_bits_manager_xact_id ),
       .io_in_6_grant_bits_is_builtin_type( outer_arb_io_in_6_grant_bits_is_builtin_type ),
       .io_in_6_grant_bits_g_type( outer_arb_io_in_6_grant_bits_g_type ),
       .io_in_6_grant_bits_data( outer_arb_io_in_6_grant_bits_data ),
       .io_in_5_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_in_5_acquire_valid( BroadcastAcquireTracker_4_io_outer_acquire_valid ),
       .io_in_5_acquire_bits_addr_block( BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_block ),
       .io_in_5_acquire_bits_client_xact_id( BroadcastAcquireTracker_4_io_outer_acquire_bits_client_xact_id ),
       .io_in_5_acquire_bits_addr_beat( BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_beat ),
       .io_in_5_acquire_bits_is_builtin_type( BroadcastAcquireTracker_4_io_outer_acquire_bits_is_builtin_type ),
       .io_in_5_acquire_bits_a_type( BroadcastAcquireTracker_4_io_outer_acquire_bits_a_type ),
       .io_in_5_acquire_bits_union( BroadcastAcquireTracker_4_io_outer_acquire_bits_union ),
       .io_in_5_acquire_bits_data( BroadcastAcquireTracker_4_io_outer_acquire_bits_data ),
       .io_in_5_grant_ready( BroadcastAcquireTracker_4_io_outer_grant_ready ),
       .io_in_5_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_in_5_grant_bits_addr_beat( outer_arb_io_in_5_grant_bits_addr_beat ),
       .io_in_5_grant_bits_client_xact_id( outer_arb_io_in_5_grant_bits_client_xact_id ),
       .io_in_5_grant_bits_manager_xact_id( outer_arb_io_in_5_grant_bits_manager_xact_id ),
       .io_in_5_grant_bits_is_builtin_type( outer_arb_io_in_5_grant_bits_is_builtin_type ),
       .io_in_5_grant_bits_g_type( outer_arb_io_in_5_grant_bits_g_type ),
       .io_in_5_grant_bits_data( outer_arb_io_in_5_grant_bits_data ),
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( BroadcastAcquireTracker_3_io_outer_acquire_valid ),
       .io_in_4_acquire_bits_addr_block( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block ),
       .io_in_4_acquire_bits_client_xact_id( BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id ),
       .io_in_4_acquire_bits_addr_beat( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat ),
       .io_in_4_acquire_bits_is_builtin_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type ),
       .io_in_4_acquire_bits_a_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type ),
       .io_in_4_acquire_bits_union( BroadcastAcquireTracker_3_io_outer_acquire_bits_union ),
       .io_in_4_acquire_bits_data( BroadcastAcquireTracker_3_io_outer_acquire_bits_data ),
       .io_in_4_grant_ready( BroadcastAcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_addr_beat( outer_arb_io_in_4_grant_bits_addr_beat ),
       .io_in_4_grant_bits_client_xact_id( outer_arb_io_in_4_grant_bits_client_xact_id ),
       .io_in_4_grant_bits_manager_xact_id( outer_arb_io_in_4_grant_bits_manager_xact_id ),
       .io_in_4_grant_bits_is_builtin_type( outer_arb_io_in_4_grant_bits_is_builtin_type ),
       .io_in_4_grant_bits_g_type( outer_arb_io_in_4_grant_bits_g_type ),
       .io_in_4_grant_bits_data( outer_arb_io_in_4_grant_bits_data ),
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( BroadcastAcquireTracker_2_io_outer_acquire_valid ),
       .io_in_3_acquire_bits_addr_block( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block ),
       .io_in_3_acquire_bits_client_xact_id( BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id ),
       .io_in_3_acquire_bits_addr_beat( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat ),
       .io_in_3_acquire_bits_is_builtin_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type ),
       .io_in_3_acquire_bits_a_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type ),
       .io_in_3_acquire_bits_union( BroadcastAcquireTracker_2_io_outer_acquire_bits_union ),
       .io_in_3_acquire_bits_data( BroadcastAcquireTracker_2_io_outer_acquire_bits_data ),
       .io_in_3_grant_ready( BroadcastAcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_addr_beat( outer_arb_io_in_3_grant_bits_addr_beat ),
       .io_in_3_grant_bits_client_xact_id( outer_arb_io_in_3_grant_bits_client_xact_id ),
       .io_in_3_grant_bits_manager_xact_id( outer_arb_io_in_3_grant_bits_manager_xact_id ),
       .io_in_3_grant_bits_is_builtin_type( outer_arb_io_in_3_grant_bits_is_builtin_type ),
       .io_in_3_grant_bits_g_type( outer_arb_io_in_3_grant_bits_g_type ),
       .io_in_3_grant_bits_data( outer_arb_io_in_3_grant_bits_data ),
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( BroadcastAcquireTracker_1_io_outer_acquire_valid ),
       .io_in_2_acquire_bits_addr_block( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block ),
       .io_in_2_acquire_bits_client_xact_id( BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id ),
       .io_in_2_acquire_bits_addr_beat( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat ),
       .io_in_2_acquire_bits_is_builtin_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type ),
       .io_in_2_acquire_bits_a_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type ),
       .io_in_2_acquire_bits_union( BroadcastAcquireTracker_1_io_outer_acquire_bits_union ),
       .io_in_2_acquire_bits_data( BroadcastAcquireTracker_1_io_outer_acquire_bits_data ),
       .io_in_2_grant_ready( BroadcastAcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_addr_beat( outer_arb_io_in_2_grant_bits_addr_beat ),
       .io_in_2_grant_bits_client_xact_id( outer_arb_io_in_2_grant_bits_client_xact_id ),
       .io_in_2_grant_bits_manager_xact_id( outer_arb_io_in_2_grant_bits_manager_xact_id ),
       .io_in_2_grant_bits_is_builtin_type( outer_arb_io_in_2_grant_bits_is_builtin_type ),
       .io_in_2_grant_bits_g_type( outer_arb_io_in_2_grant_bits_g_type ),
       .io_in_2_grant_bits_data( outer_arb_io_in_2_grant_bits_data ),
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( BroadcastAcquireTracker_io_outer_acquire_valid ),
       .io_in_1_acquire_bits_addr_block( BroadcastAcquireTracker_io_outer_acquire_bits_addr_block ),
       .io_in_1_acquire_bits_client_xact_id( BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id ),
       .io_in_1_acquire_bits_addr_beat( BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat ),
       .io_in_1_acquire_bits_is_builtin_type( BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_in_1_acquire_bits_a_type( BroadcastAcquireTracker_io_outer_acquire_bits_a_type ),
       .io_in_1_acquire_bits_union( BroadcastAcquireTracker_io_outer_acquire_bits_union ),
       .io_in_1_acquire_bits_data( BroadcastAcquireTracker_io_outer_acquire_bits_data ),
       .io_in_1_grant_ready( BroadcastAcquireTracker_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_addr_beat( outer_arb_io_in_1_grant_bits_addr_beat ),
       .io_in_1_grant_bits_client_xact_id( outer_arb_io_in_1_grant_bits_client_xact_id ),
       .io_in_1_grant_bits_manager_xact_id( outer_arb_io_in_1_grant_bits_manager_xact_id ),
       .io_in_1_grant_bits_is_builtin_type( outer_arb_io_in_1_grant_bits_is_builtin_type ),
       .io_in_1_grant_bits_g_type( outer_arb_io_in_1_grant_bits_g_type ),
       .io_in_1_grant_bits_data( outer_arb_io_in_1_grant_bits_data ),
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_in_0_acquire_bits_addr_block( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block ),
       .io_in_0_acquire_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id ),
       .io_in_0_acquire_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat ),
       .io_in_0_acquire_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_in_0_acquire_bits_a_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type ),
       .io_in_0_acquire_bits_union( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union ),
       .io_in_0_acquire_bits_data( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data ),
       .io_in_0_grant_ready( BroadcastVoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_addr_beat( outer_arb_io_in_0_grant_bits_addr_beat ),
       .io_in_0_grant_bits_client_xact_id( outer_arb_io_in_0_grant_bits_client_xact_id ),
       .io_in_0_grant_bits_manager_xact_id( outer_arb_io_in_0_grant_bits_manager_xact_id ),
       .io_in_0_grant_bits_is_builtin_type( outer_arb_io_in_0_grant_bits_is_builtin_type ),
       .io_in_0_grant_bits_g_type( outer_arb_io_in_0_grant_bits_g_type ),
       .io_in_0_grant_bits_data( outer_arb_io_in_0_grant_bits_data ),
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( outer_arb_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( outer_arb_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( outer_arb_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( outer_arb_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( outer_arb_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( outer_arb_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( outer_arb_io_out_acquire_bits_data ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_addr_beat( io_outer_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( io_outer_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( io_outer_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( io_outer_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( io_outer_grant_bits_g_type ),
       .io_out_grant_bits_data( T293 )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Non-voluntary release should always have a Tracker waiting for it.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      rel_data_cnt <= 2'h0;
    end else if(vwbdq_enq) begin
      rel_data_cnt <= T18;
    end
    if(reset) begin
      sdq_val <= 4'h0;
    end else if(T72) begin
      sdq_val <= T36;
    end
    if(T221) begin
      vwbdq_0 <= io_inner_release_bits_data;
    end
    if(T226) begin
      vwbdq_1 <= io_inner_release_bits_data;
    end
    if(T232) begin
      vwbdq_2 <= io_inner_release_bits_data;
    end
    if(T235) begin
      vwbdq_3 <= io_inner_release_bits_data;
    end
    if(T243) begin
      sdq_0 <= io_inner_acquire_bits_data;
    end
    if(T248) begin
      sdq_1 <= io_inner_acquire_bits_data;
    end
    if(T254) begin
      sdq_2 <= io_inner_acquire_bits_data;
    end
    if(T257) begin
      sdq_3 <= io_inner_acquire_bits_data;
    end
  end
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [31:0] io_enq_bits_addr,
    input [7:0] io_enq_bits_len,
    input [2:0] io_enq_bits_size,
    input [1:0] io_enq_bits_burst,
    input  io_enq_bits_lock,
    input [3:0] io_enq_bits_cache,
    input [2:0] io_enq_bits_prot,
    input [3:0] io_enq_bits_qos,
    input [3:0] io_enq_bits_region,
    input [4:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[31:0] io_deq_bits_addr,
    output[7:0] io_deq_bits_len,
    output[2:0] io_deq_bits_size,
    output[1:0] io_deq_bits_burst,
    output io_deq_bits_lock,
    output[3:0] io_deq_bits_cache,
    output[2:0] io_deq_bits_prot,
    output[3:0] io_deq_bits_qos,
    output[3:0] io_deq_bits_region,
    output[4:0] io_deq_bits_id,
    output io_deq_bits_user,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T37;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T38;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T39;
  wire T8;
  wire T9;
  wire T10;
  wire[66:0] T11;
  reg [66:0] ram [1:0];
  wire[66:0] T12;
  wire[66:0] T13;
  wire[66:0] T14;
  wire[20:0] T15;
  wire[9:0] T16;
  wire[5:0] T17;
  wire[10:0] T18;
  wire[6:0] T19;
  wire[45:0] T20;
  wire[5:0] T21;
  wire[2:0] T22;
  wire[39:0] T23;
  wire[4:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[2:0] T27;
  wire[3:0] T28;
  wire T29;
  wire[1:0] T30;
  wire[2:0] T31;
  wire[7:0] T32;
  wire[31:0] T33;
  wire T34;
  wire empty;
  wire T35;
  wire T36;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T37 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T38 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T39 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T20, T15};
  assign T15 = {T18, T16};
  assign T16 = {io_enq_bits_region, T17};
  assign T17 = {io_enq_bits_id, io_enq_bits_user};
  assign T18 = {io_enq_bits_cache, T19};
  assign T19 = {io_enq_bits_prot, io_enq_bits_qos};
  assign T20 = {T23, T21};
  assign T21 = {io_enq_bits_size, T22};
  assign T22 = {io_enq_bits_burst, io_enq_bits_lock};
  assign T23 = {io_enq_bits_addr, io_enq_bits_len};
  assign io_deq_bits_id = T24;
  assign T24 = T11[3'h5:1'h1];
  assign io_deq_bits_region = T25;
  assign T25 = T11[4'h9:3'h6];
  assign io_deq_bits_qos = T26;
  assign T26 = T11[4'hd:4'ha];
  assign io_deq_bits_prot = T27;
  assign T27 = T11[5'h10:4'he];
  assign io_deq_bits_cache = T28;
  assign T28 = T11[5'h14:5'h11];
  assign io_deq_bits_lock = T29;
  assign T29 = T11[5'h15:5'h15];
  assign io_deq_bits_burst = T30;
  assign T30 = T11[5'h17:5'h16];
  assign io_deq_bits_size = T31;
  assign T31 = T11[5'h1a:5'h18];
  assign io_deq_bits_len = T32;
  assign T32 = T11[6'h22:5'h1b];
  assign io_deq_bits_addr = T33;
  assign T33 = T11[7'h42:6'h23];
  assign io_deq_valid = T34;
  assign T34 = empty ^ 1'h1;
  assign empty = ptr_match & T35;
  assign T35 = maybe_full ^ 1'h1;
  assign io_enq_ready = T36;
  assign T36 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [4:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[4:0] io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire[4:0] T10;
  reg [4:0] ram [1:0];
  wire[4:0] T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module NastiErrorSlave(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [4:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    output[1:0] io_b_bits_resp,
    output[4:0] io_b_bits_id,
    //output io_b_bits_user
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [4:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[4:0] io_r_bits_id
    //output io_r_bits_user
);

  wire T0;
  wire T1;
  wire T2;
  wire[31:0] T3;
  wire[247:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire[31:0] T8;
  wire[239:0] T9;
  wire T10;
  wire T11;
  reg  draining;
  wire T39;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  reg [7:0] beats_left;
  wire[7:0] T40;
  wire[7:0] T22;
  wire[7:0] T23;
  wire T24;
  wire T25;
  reg  responding;
  wire T41;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire r_queue_io_enq_ready;
  wire r_queue_io_deq_valid;
  wire[7:0] r_queue_io_deq_bits_len;
  wire[4:0] r_queue_io_deq_bits_id;
  wire b_queue_io_enq_ready;
  wire b_queue_io_deq_valid;
  wire[4:0] b_queue_io_deq_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    draining = {1{$random}};
    beats_left = {1{$random}};
    responding = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_r_bits_user = {1{$random}};
//  assign io_b_bits_user = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T2 & T1;
  assign T1 = reset ^ 1'h1;
  assign T2 = io_aw_ready & io_aw_valid;
  assign T3 = io_aw_bits_addr;
  assign T5 = T7 & T6;
  assign T6 = reset ^ 1'h1;
  assign T7 = io_ar_ready & io_ar_valid;
  assign T8 = io_ar_bits_addr;
  assign T10 = io_b_ready & T11;
  assign T11 = draining ^ 1'h1;
  assign T39 = reset ? 1'h0 : T12;
  assign T12 = T15 ? 1'h0 : T13;
  assign T13 = T14 ? 1'h1 : draining;
  assign T14 = io_aw_ready & io_aw_valid;
  assign T15 = T16 & io_w_bits_last;
  assign T16 = io_w_ready & io_w_valid;
  assign T17 = io_aw_valid & T18;
  assign T18 = draining ^ 1'h1;
  assign T19 = T20 & io_r_bits_last;
  assign T20 = io_r_ready & io_r_valid;
  assign io_r_bits_id = r_queue_io_deq_bits_id;
  assign io_r_bits_last = T21;
  assign T21 = beats_left == 8'h0;
  assign T40 = reset ? 8'h0 : T22;
  assign T22 = T32 ? T31 : T23;
  assign T23 = T24 ? r_queue_io_deq_bits_len : beats_left;
  assign T24 = T25 & r_queue_io_deq_valid;
  assign T25 = responding ^ 1'h1;
  assign T41 = reset ? 1'h0 : T26;
  assign T26 = T28 ? 1'h0 : T27;
  assign T27 = T24 ? 1'h1 : responding;
  assign T28 = T30 & T29;
  assign T29 = beats_left == 8'h0;
  assign T30 = io_r_ready & io_r_valid;
  assign T31 = beats_left - 8'h0;
  assign T32 = T30 & T33;
  assign T33 = T29 ^ 1'h1;
  assign io_r_bits_data = 64'h0;
  assign io_r_bits_resp = 2'h3;
  assign io_r_valid = T34;
  assign T34 = r_queue_io_deq_valid & responding;
  assign io_ar_ready = r_queue_io_enq_ready;
  assign io_b_bits_id = b_queue_io_deq_bits;
  assign io_b_bits_resp = 2'h3;
  assign io_b_valid = T35;
  assign T35 = b_queue_io_deq_valid & T36;
  assign T36 = draining ^ 1'h1;
  assign io_w_ready = draining;
  assign io_aw_ready = T37;
  assign T37 = b_queue_io_enq_ready & T38;
  assign T38 = draining ^ 1'h1;
  Queue_3 r_queue(.clk(clk), .reset(reset),
       .io_enq_ready( r_queue_io_enq_ready ),
       .io_enq_valid( io_ar_valid ),
       .io_enq_bits_addr( io_ar_bits_addr ),
       .io_enq_bits_len( io_ar_bits_len ),
       .io_enq_bits_size( io_ar_bits_size ),
       .io_enq_bits_burst( io_ar_bits_burst ),
       .io_enq_bits_lock( io_ar_bits_lock ),
       .io_enq_bits_cache( io_ar_bits_cache ),
       .io_enq_bits_prot( io_ar_bits_prot ),
       .io_enq_bits_qos( io_ar_bits_qos ),
       .io_enq_bits_region( io_ar_bits_region ),
       .io_enq_bits_id( io_ar_bits_id ),
       .io_enq_bits_user( io_ar_bits_user ),
       .io_deq_ready( T19 ),
       .io_deq_valid( r_queue_io_deq_valid ),
       //.io_deq_bits_addr(  )
       .io_deq_bits_len( r_queue_io_deq_bits_len ),
       //.io_deq_bits_size(  )
       //.io_deq_bits_burst(  )
       //.io_deq_bits_lock(  )
       //.io_deq_bits_cache(  )
       //.io_deq_bits_prot(  )
       //.io_deq_bits_qos(  )
       //.io_deq_bits_region(  )
       .io_deq_bits_id( r_queue_io_deq_bits_id )
       //.io_deq_bits_user(  )
       //.io_count(  )
  );
  Queue_7 b_queue(.clk(clk), .reset(reset),
       .io_enq_ready( b_queue_io_enq_ready ),
       .io_enq_valid( T17 ),
       .io_enq_bits( io_aw_bits_id ),
       .io_deq_ready( T10 ),
       .io_deq_valid( b_queue_io_deq_valid ),
       .io_deq_bits( b_queue_io_deq_bits )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      draining <= 1'h0;
    end else if(T15) begin
      draining <= 1'h0;
    end else if(T14) begin
      draining <= 1'h1;
    end
    if(reset) begin
      beats_left <= 8'h0;
    end else if(T32) begin
      beats_left <= T31;
    end else if(T24) begin
      beats_left <= r_queue_io_deq_bits_len;
    end
    if(reset) begin
      responding <= 1'h0;
    end else if(T28) begin
      responding <= 1'h0;
    end else if(T24) begin
      responding <= 1'h1;
    end
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T5)
        $fwrite(32'h80000002, "Invalid read address %h\n", T8);
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "Invalid write address %h\n", T3);
// synthesis translate_on
`endif
  end
endmodule

module RRArbiter_4(input clk, input reset,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_resp,
    input [4:0] io_in_3_bits_id,
    input  io_in_3_bits_user,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [4:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [4:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [4:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[4:0] io_out_bits_id,
    output io_out_bits_user,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg [1:0] last_grant;
  wire[1:0] T89;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[4:0] T20;
  wire[4:0] T21;
  wire T22;
  wire[4:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T11 ? 2'h1 : T0;
  assign T0 = T9 ? 2'h2 : T1;
  assign T1 = T5 ? 2'h3 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : T4;
  assign T4 = io_in_2_valid ? 2'h2 : 2'h3;
  assign T5 = io_in_3_valid & T6;
  assign T6 = last_grant < 2'h3;
  assign T89 = reset ? 2'h0 : T7;
  assign T7 = T8 ? chosen : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_2_valid & T10;
  assign T10 = last_grant < 2'h2;
  assign T11 = io_in_1_valid & T12;
  assign T12 = last_grant < 2'h1;
  assign io_out_bits_user = T13;
  assign T13 = T19 ? T17 : T14;
  assign T14 = T15 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T15 = T16[1'h0:1'h0];
  assign T16 = chosen;
  assign T17 = T18 ? io_in_3_bits_user : io_in_2_bits_user;
  assign T18 = T16[1'h0:1'h0];
  assign T19 = T16[1'h1:1'h1];
  assign io_out_bits_id = T20;
  assign T20 = T25 ? T23 : T21;
  assign T21 = T22 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T22 = T16[1'h0:1'h0];
  assign T23 = T24 ? io_in_3_bits_id : io_in_2_bits_id;
  assign T24 = T16[1'h0:1'h0];
  assign T25 = T16[1'h1:1'h1];
  assign io_out_bits_resp = T26;
  assign T26 = T31 ? T29 : T27;
  assign T27 = T28 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T28 = T16[1'h0:1'h0];
  assign T29 = T30 ? io_in_3_bits_resp : io_in_2_bits_resp;
  assign T30 = T16[1'h0:1'h0];
  assign T31 = T16[1'h1:1'h1];
  assign io_out_valid = T32;
  assign T32 = T37 ? T35 : T33;
  assign T33 = T34 ? io_in_1_valid : io_in_0_valid;
  assign T34 = T16[1'h0:1'h0];
  assign T35 = T36 ? io_in_3_valid : io_in_2_valid;
  assign T36 = T16[1'h0:1'h0];
  assign T37 = T16[1'h1:1'h1];
  assign io_in_0_ready = T38;
  assign T38 = T39 & io_out_ready;
  assign T39 = T52 | T40;
  assign T40 = T41 ^ 1'h1;
  assign T41 = T44 | T42;
  assign T42 = io_in_3_valid & T43;
  assign T43 = last_grant < 2'h3;
  assign T44 = T47 | T45;
  assign T45 = io_in_2_valid & T46;
  assign T46 = last_grant < 2'h2;
  assign T47 = T50 | T48;
  assign T48 = io_in_1_valid & T49;
  assign T49 = last_grant < 2'h1;
  assign T50 = io_in_0_valid & T51;
  assign T51 = last_grant < 2'h0;
  assign T52 = last_grant < 2'h0;
  assign io_in_1_ready = T53;
  assign T53 = T54 & io_out_ready;
  assign T54 = T60 | T55;
  assign T55 = T56 ^ 1'h1;
  assign T56 = T57 | io_in_0_valid;
  assign T57 = T58 | T42;
  assign T58 = T59 | T45;
  assign T59 = T50 | T48;
  assign T60 = T62 & T61;
  assign T61 = last_grant < 2'h1;
  assign T62 = T50 ^ 1'h1;
  assign io_in_2_ready = T63;
  assign T63 = T64 & io_out_ready;
  assign T64 = T71 | T65;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_1_valid;
  assign T67 = T68 | io_in_0_valid;
  assign T68 = T69 | T42;
  assign T69 = T70 | T45;
  assign T70 = T50 | T48;
  assign T71 = T73 & T72;
  assign T72 = last_grant < 2'h2;
  assign T73 = T74 ^ 1'h1;
  assign T74 = T50 | T48;
  assign io_in_3_ready = T75;
  assign T75 = T76 & io_out_ready;
  assign T76 = T84 | T77;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T79 | io_in_2_valid;
  assign T79 = T80 | io_in_1_valid;
  assign T80 = T81 | io_in_0_valid;
  assign T81 = T82 | T42;
  assign T82 = T83 | T45;
  assign T83 = T50 | T48;
  assign T84 = T86 & T85;
  assign T85 = last_grant < 2'h3;
  assign T86 = T87 ^ 1'h1;
  assign T87 = T88 | T45;
  assign T88 = T50 | T48;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= chosen;
    end
  end
endmodule

module JunctionsPeekingArbiter_0(input clk, input reset,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_resp,
    input [63:0] io_in_3_bits_data,
    input  io_in_3_bits_last,
    input [4:0] io_in_3_bits_id,
    input  io_in_3_bits_user,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [63:0] io_in_2_bits_data,
    input  io_in_2_bits_last,
    input [4:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [63:0] io_in_1_bits_data,
    input  io_in_1_bits_last,
    input [4:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_last,
    input [4:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[63:0] io_out_bits_data,
    output io_out_bits_last,
    output[4:0] io_out_bits_id,
    output io_out_bits_user
);

  wire T0;
  wire T1;
  wire T2;
  wire[1:0] T3;
  wire[1:0] chosen;
  wire[1:0] choice;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  reg [1:0] T7;
  wire[1:0] T9;
  wire[1:0] T10;
  reg [1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  reg [1:0] T15;
  wire[1:0] T16;
  reg [1:0] T17;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  reg [1:0] T40;
  wire[1:0] T41;
  reg [1:0] T42;
  wire[1:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[1:0] T63;
  reg [1:0] T64;
  wire[1:0] T135;
  wire[2:0] T65;
  wire[2:0] T136;
  reg [1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[2:0] T137;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[1:0] T73;
  wire[1:0] T138;
  wire[2:0] T74;
  wire[2:0] T139;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[2:0] T140;
  reg [1:0] lockIdx;
  wire[1:0] T141;
  wire[1:0] T87;
  wire T88;
  wire T89;
  wire T90;
  reg  locked;
  wire T142;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire[4:0] T97;
  wire[4:0] T98;
  wire T99;
  wire[4:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[63:0] T109;
  wire[63:0] T110;
  wire T111;
  wire[63:0] T112;
  wire T113;
  wire T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_bits_user = T0;
  assign T0 = T96 ? T94 : T1;
  assign T1 = T2 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T2 = T3[1'h0:1'h0];
  assign T3 = chosen;
  assign chosen = locked ? lockIdx : choice;
  assign choice = T69 ? T63 : T4;
  assign T4 = T45 ? T39 : T5;
  assign T5 = T20 ? T14 : T6;
  assign T6 = T13 ? T11 : T7;
  always @(*) case (T9)
    0: T7 = 2'h0;
    1: T7 = 2'h1;
    2: T7 = 2'h2;
    3: T7 = 2'h3;
    default: begin
      T7 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T7 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T9 = T10 - 2'h1;
  assign T10 = lockIdx + 2'h1;
  always @(*) case (T12)
    0: T11 = 2'h0;
    1: T11 = 2'h1;
    2: T11 = 2'h2;
    3: T11 = 2'h3;
    default: begin
      T11 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T11 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T12 = 2'h3 + T10;
  assign T13 = T10 < 2'h1;
  assign T14 = T19 ? T17 : T15;
  always @(*) case (T16)
    0: T15 = 2'h0;
    1: T15 = 2'h1;
    2: T15 = 2'h2;
    3: T15 = 2'h3;
    default: begin
      T15 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T15 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T16 = T10 - 2'h2;
  always @(*) case (T18)
    0: T17 = 2'h0;
    1: T17 = 2'h1;
    2: T17 = 2'h2;
    3: T17 = 2'h3;
    default: begin
      T17 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T17 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T18 = 2'h2 + T10;
  assign T19 = T10 < 2'h2;
  assign T20 = T38 ? T30 : T21;
  assign T21 = T29 ? T27 : T22;
  assign T22 = T23 ? io_in_1_valid : io_in_0_valid;
  assign T23 = T24[1'h0:1'h0];
  assign T24 = T25;
  assign T25 = T26 - 2'h2;
  assign T26 = lockIdx + 2'h1;
  assign T27 = T28 ? io_in_3_valid : io_in_2_valid;
  assign T28 = T24[1'h0:1'h0];
  assign T29 = T24[1'h1:1'h1];
  assign T30 = T37 ? T35 : T31;
  assign T31 = T32 ? io_in_1_valid : io_in_0_valid;
  assign T32 = T33[1'h0:1'h0];
  assign T33 = T34;
  assign T34 = 2'h2 + T26;
  assign T35 = T36 ? io_in_3_valid : io_in_2_valid;
  assign T36 = T33[1'h0:1'h0];
  assign T37 = T33[1'h1:1'h1];
  assign T38 = T26 < 2'h2;
  assign T39 = T44 ? T42 : T40;
  always @(*) case (T41)
    0: T40 = 2'h0;
    1: T40 = 2'h1;
    2: T40 = 2'h2;
    3: T40 = 2'h3;
    default: begin
      T40 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T40 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T41 = T10 - 2'h3;
  always @(*) case (T43)
    0: T42 = 2'h0;
    1: T42 = 2'h1;
    2: T42 = 2'h2;
    3: T42 = 2'h3;
    default: begin
      T42 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T42 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T43 = 2'h1 + T10;
  assign T44 = T10 < 2'h3;
  assign T45 = T62 ? T54 : T46;
  assign T46 = T53 ? T51 : T47;
  assign T47 = T48 ? io_in_1_valid : io_in_0_valid;
  assign T48 = T49[1'h0:1'h0];
  assign T49 = T50;
  assign T50 = T26 - 2'h3;
  assign T51 = T52 ? io_in_3_valid : io_in_2_valid;
  assign T52 = T49[1'h0:1'h0];
  assign T53 = T49[1'h1:1'h1];
  assign T54 = T61 ? T59 : T55;
  assign T55 = T56 ? io_in_1_valid : io_in_0_valid;
  assign T56 = T57[1'h0:1'h0];
  assign T57 = T58;
  assign T58 = 2'h1 + T26;
  assign T59 = T60 ? io_in_3_valid : io_in_2_valid;
  assign T60 = T57[1'h0:1'h0];
  assign T61 = T57[1'h1:1'h1];
  assign T62 = T26 < 2'h3;
  assign T63 = T68 ? T66 : T64;
  always @(*) case (T135)
    0: T64 = 2'h0;
    1: T64 = 2'h1;
    2: T64 = 2'h2;
    3: T64 = 2'h3;
    default: begin
      T64 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T64 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T135 = T65[1'h1:1'h0];
  assign T65 = T136 - 3'h4;
  assign T136 = {1'h0, T10};
  always @(*) case (T67)
    0: T66 = 2'h0;
    1: T66 = 2'h1;
    2: T66 = 2'h2;
    3: T66 = 2'h3;
    default: begin
      T66 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T66 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T67 = 2'h0 + T10;
  assign T68 = T137 < 3'h4;
  assign T137 = {1'h0, T10};
  assign T69 = T86 ? T78 : T70;
  assign T70 = T77 ? T75 : T71;
  assign T71 = T72 ? io_in_1_valid : io_in_0_valid;
  assign T72 = T73[1'h0:1'h0];
  assign T73 = T138;
  assign T138 = T74[1'h1:1'h0];
  assign T74 = T139 - 3'h4;
  assign T139 = {1'h0, T26};
  assign T75 = T76 ? io_in_3_valid : io_in_2_valid;
  assign T76 = T73[1'h0:1'h0];
  assign T77 = T73[1'h1:1'h1];
  assign T78 = T85 ? T83 : T79;
  assign T79 = T80 ? io_in_1_valid : io_in_0_valid;
  assign T80 = T81[1'h0:1'h0];
  assign T81 = T82;
  assign T82 = 2'h0 + T26;
  assign T83 = T84 ? io_in_3_valid : io_in_2_valid;
  assign T84 = T81[1'h0:1'h0];
  assign T85 = T81[1'h1:1'h1];
  assign T86 = T140 < 3'h4;
  assign T140 = {1'h0, T26};
  assign T141 = reset ? 2'h0 : T87;
  assign T87 = T88 ? choice : lockIdx;
  assign T88 = T90 & T89;
  assign T89 = locked ^ 1'h1;
  assign T90 = io_out_ready & io_out_valid;
  assign T142 = reset ? 1'h0 : T91;
  assign T91 = T93 ? 1'h0 : T92;
  assign T92 = T88 ? 1'h1 : locked;
  assign T93 = T90 & io_out_bits_last;
  assign T94 = T95 ? io_in_3_bits_user : io_in_2_bits_user;
  assign T95 = T3[1'h0:1'h0];
  assign T96 = T3[1'h1:1'h1];
  assign io_out_bits_id = T97;
  assign T97 = T102 ? T100 : T98;
  assign T98 = T99 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T99 = T3[1'h0:1'h0];
  assign T100 = T101 ? io_in_3_bits_id : io_in_2_bits_id;
  assign T101 = T3[1'h0:1'h0];
  assign T102 = T3[1'h1:1'h1];
  assign io_out_bits_last = T103;
  assign T103 = T108 ? T106 : T104;
  assign T104 = T105 ? io_in_1_bits_last : io_in_0_bits_last;
  assign T105 = T3[1'h0:1'h0];
  assign T106 = T107 ? io_in_3_bits_last : io_in_2_bits_last;
  assign T107 = T3[1'h0:1'h0];
  assign T108 = T3[1'h1:1'h1];
  assign io_out_bits_data = T109;
  assign T109 = T114 ? T112 : T110;
  assign T110 = T111 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T111 = T3[1'h0:1'h0];
  assign T112 = T113 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T113 = T3[1'h0:1'h0];
  assign T114 = T3[1'h1:1'h1];
  assign io_out_bits_resp = T115;
  assign T115 = T120 ? T118 : T116;
  assign T116 = T117 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T117 = T3[1'h0:1'h0];
  assign T118 = T119 ? io_in_3_bits_resp : io_in_2_bits_resp;
  assign T119 = T3[1'h0:1'h0];
  assign T120 = T3[1'h1:1'h1];
  assign io_out_valid = T121;
  assign T121 = T126 ? T124 : T122;
  assign T122 = T123 ? io_in_1_valid : io_in_0_valid;
  assign T123 = T3[1'h0:1'h0];
  assign T124 = T125 ? io_in_3_valid : io_in_2_valid;
  assign T125 = T3[1'h0:1'h0];
  assign T126 = T3[1'h1:1'h1];
  assign io_in_0_ready = T127;
  assign T127 = io_out_ready & T128;
  assign T128 = chosen == 2'h0;
  assign io_in_1_ready = T129;
  assign T129 = io_out_ready & T130;
  assign T130 = chosen == 2'h1;
  assign io_in_2_ready = T131;
  assign T131 = io_out_ready & T132;
  assign T132 = chosen == 2'h2;
  assign io_in_3_ready = T133;
  assign T133 = io_out_ready & T134;
  assign T134 = chosen == 2'h3;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 2'h0;
    end else if(T88) begin
      lockIdx <= choice;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T93) begin
      locked <= 1'h0;
    end else if(T88) begin
      locked <= 1'h1;
    end
  end
endmodule

module NastiRouter_0(input clk, input reset,
    output io_master_aw_ready,
    input  io_master_aw_valid,
    input [31:0] io_master_aw_bits_addr,
    input [7:0] io_master_aw_bits_len,
    input [2:0] io_master_aw_bits_size,
    input [1:0] io_master_aw_bits_burst,
    input  io_master_aw_bits_lock,
    input [3:0] io_master_aw_bits_cache,
    input [2:0] io_master_aw_bits_prot,
    input [3:0] io_master_aw_bits_qos,
    input [3:0] io_master_aw_bits_region,
    input [4:0] io_master_aw_bits_id,
    input  io_master_aw_bits_user,
    output io_master_w_ready,
    input  io_master_w_valid,
    input [63:0] io_master_w_bits_data,
    input  io_master_w_bits_last,
    input [7:0] io_master_w_bits_strb,
    input  io_master_w_bits_user,
    input  io_master_b_ready,
    output io_master_b_valid,
    output[1:0] io_master_b_bits_resp,
    output[4:0] io_master_b_bits_id,
    output io_master_b_bits_user,
    output io_master_ar_ready,
    input  io_master_ar_valid,
    input [31:0] io_master_ar_bits_addr,
    input [7:0] io_master_ar_bits_len,
    input [2:0] io_master_ar_bits_size,
    input [1:0] io_master_ar_bits_burst,
    input  io_master_ar_bits_lock,
    input [3:0] io_master_ar_bits_cache,
    input [2:0] io_master_ar_bits_prot,
    input [3:0] io_master_ar_bits_qos,
    input [3:0] io_master_ar_bits_region,
    input [4:0] io_master_ar_bits_id,
    input  io_master_ar_bits_user,
    input  io_master_r_ready,
    output io_master_r_valid,
    output[1:0] io_master_r_bits_resp,
    output[63:0] io_master_r_bits_data,
    output io_master_r_bits_last,
    output[4:0] io_master_r_bits_id,
    output io_master_r_bits_user,
    input  io_slave_2_aw_ready,
    output io_slave_2_aw_valid,
    output[31:0] io_slave_2_aw_bits_addr,
    output[7:0] io_slave_2_aw_bits_len,
    output[2:0] io_slave_2_aw_bits_size,
    output[1:0] io_slave_2_aw_bits_burst,
    output io_slave_2_aw_bits_lock,
    output[3:0] io_slave_2_aw_bits_cache,
    output[2:0] io_slave_2_aw_bits_prot,
    output[3:0] io_slave_2_aw_bits_qos,
    output[3:0] io_slave_2_aw_bits_region,
    output[4:0] io_slave_2_aw_bits_id,
    output io_slave_2_aw_bits_user,
    input  io_slave_2_w_ready,
    output io_slave_2_w_valid,
    output[63:0] io_slave_2_w_bits_data,
    output io_slave_2_w_bits_last,
    output[7:0] io_slave_2_w_bits_strb,
    output io_slave_2_w_bits_user,
    output io_slave_2_b_ready,
    input  io_slave_2_b_valid,
    input [1:0] io_slave_2_b_bits_resp,
    input [4:0] io_slave_2_b_bits_id,
    input  io_slave_2_b_bits_user,
    input  io_slave_2_ar_ready,
    output io_slave_2_ar_valid,
    output[31:0] io_slave_2_ar_bits_addr,
    output[7:0] io_slave_2_ar_bits_len,
    output[2:0] io_slave_2_ar_bits_size,
    output[1:0] io_slave_2_ar_bits_burst,
    output io_slave_2_ar_bits_lock,
    output[3:0] io_slave_2_ar_bits_cache,
    output[2:0] io_slave_2_ar_bits_prot,
    output[3:0] io_slave_2_ar_bits_qos,
    output[3:0] io_slave_2_ar_bits_region,
    output[4:0] io_slave_2_ar_bits_id,
    output io_slave_2_ar_bits_user,
    output io_slave_2_r_ready,
    input  io_slave_2_r_valid,
    input [1:0] io_slave_2_r_bits_resp,
    input [63:0] io_slave_2_r_bits_data,
    input  io_slave_2_r_bits_last,
    input [4:0] io_slave_2_r_bits_id,
    input  io_slave_2_r_bits_user,
    input  io_slave_1_aw_ready,
    output io_slave_1_aw_valid,
    output[31:0] io_slave_1_aw_bits_addr,
    output[7:0] io_slave_1_aw_bits_len,
    output[2:0] io_slave_1_aw_bits_size,
    output[1:0] io_slave_1_aw_bits_burst,
    output io_slave_1_aw_bits_lock,
    output[3:0] io_slave_1_aw_bits_cache,
    output[2:0] io_slave_1_aw_bits_prot,
    output[3:0] io_slave_1_aw_bits_qos,
    output[3:0] io_slave_1_aw_bits_region,
    output[4:0] io_slave_1_aw_bits_id,
    output io_slave_1_aw_bits_user,
    input  io_slave_1_w_ready,
    output io_slave_1_w_valid,
    output[63:0] io_slave_1_w_bits_data,
    output io_slave_1_w_bits_last,
    output[7:0] io_slave_1_w_bits_strb,
    output io_slave_1_w_bits_user,
    output io_slave_1_b_ready,
    input  io_slave_1_b_valid,
    input [1:0] io_slave_1_b_bits_resp,
    input [4:0] io_slave_1_b_bits_id,
    input  io_slave_1_b_bits_user,
    input  io_slave_1_ar_ready,
    output io_slave_1_ar_valid,
    output[31:0] io_slave_1_ar_bits_addr,
    output[7:0] io_slave_1_ar_bits_len,
    output[2:0] io_slave_1_ar_bits_size,
    output[1:0] io_slave_1_ar_bits_burst,
    output io_slave_1_ar_bits_lock,
    output[3:0] io_slave_1_ar_bits_cache,
    output[2:0] io_slave_1_ar_bits_prot,
    output[3:0] io_slave_1_ar_bits_qos,
    output[3:0] io_slave_1_ar_bits_region,
    output[4:0] io_slave_1_ar_bits_id,
    output io_slave_1_ar_bits_user,
    output io_slave_1_r_ready,
    input  io_slave_1_r_valid,
    input [1:0] io_slave_1_r_bits_resp,
    input [63:0] io_slave_1_r_bits_data,
    input  io_slave_1_r_bits_last,
    input [4:0] io_slave_1_r_bits_id,
    input  io_slave_1_r_bits_user,
    input  io_slave_0_aw_ready,
    output io_slave_0_aw_valid,
    output[31:0] io_slave_0_aw_bits_addr,
    output[7:0] io_slave_0_aw_bits_len,
    output[2:0] io_slave_0_aw_bits_size,
    output[1:0] io_slave_0_aw_bits_burst,
    output io_slave_0_aw_bits_lock,
    output[3:0] io_slave_0_aw_bits_cache,
    output[2:0] io_slave_0_aw_bits_prot,
    output[3:0] io_slave_0_aw_bits_qos,
    output[3:0] io_slave_0_aw_bits_region,
    output[4:0] io_slave_0_aw_bits_id,
    output io_slave_0_aw_bits_user,
    input  io_slave_0_w_ready,
    output io_slave_0_w_valid,
    output[63:0] io_slave_0_w_bits_data,
    output io_slave_0_w_bits_last,
    output[7:0] io_slave_0_w_bits_strb,
    output io_slave_0_w_bits_user,
    output io_slave_0_b_ready,
    input  io_slave_0_b_valid,
    input [1:0] io_slave_0_b_bits_resp,
    input [4:0] io_slave_0_b_bits_id,
    input  io_slave_0_b_bits_user,
    input  io_slave_0_ar_ready,
    output io_slave_0_ar_valid,
    output[31:0] io_slave_0_ar_bits_addr,
    output[7:0] io_slave_0_ar_bits_len,
    output[2:0] io_slave_0_ar_bits_size,
    output[1:0] io_slave_0_ar_bits_burst,
    output io_slave_0_ar_bits_lock,
    output[3:0] io_slave_0_ar_bits_cache,
    output[2:0] io_slave_0_ar_bits_prot,
    output[3:0] io_slave_0_ar_bits_qos,
    output[3:0] io_slave_0_ar_bits_region,
    output[4:0] io_slave_0_ar_bits_id,
    output io_slave_0_ar_bits_user,
    output io_slave_0_r_ready,
    input  io_slave_0_r_valid,
    input [1:0] io_slave_0_r_bits_resp,
    input [63:0] io_slave_0_r_bits_data,
    input  io_slave_0_r_bits_last,
    input [4:0] io_slave_0_r_bits_id,
    input  io_slave_0_r_bits_user
);

  wire T0;
  wire r_invalid;
  wire T1;
  wire[2:0] ar_route;
  wire[2:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[32:0] T82;
  wire T12;
  wire T13;
  wire w_invalid;
  wire T14;
  wire[2:0] aw_route;
  wire[2:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[32:0] T83;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  reg  R29;
  wire T84;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  reg  R40;
  wire T85;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  reg  R51;
  wire T86;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire ar_ready;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire w_ready;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire aw_ready;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire b_arb_io_in_3_ready;
  wire b_arb_io_in_2_ready;
  wire b_arb_io_in_1_ready;
  wire b_arb_io_in_0_ready;
  wire b_arb_io_out_valid;
  wire[1:0] b_arb_io_out_bits_resp;
  wire[4:0] b_arb_io_out_bits_id;
  wire b_arb_io_out_bits_user;
  wire r_arb_io_in_3_ready;
  wire r_arb_io_in_2_ready;
  wire r_arb_io_in_1_ready;
  wire r_arb_io_in_0_ready;
  wire r_arb_io_out_valid;
  wire[1:0] r_arb_io_out_bits_resp;
  wire[63:0] r_arb_io_out_bits_data;
  wire r_arb_io_out_bits_last;
  wire[4:0] r_arb_io_out_bits_id;
  wire r_arb_io_out_bits_user;
  wire err_slave_io_aw_ready;
  wire err_slave_io_w_ready;
  wire err_slave_io_b_valid;
  wire[1:0] err_slave_io_b_bits_resp;
  wire[4:0] err_slave_io_b_bits_id;
  wire err_slave_io_ar_ready;
  wire err_slave_io_r_valid;
  wire[1:0] err_slave_io_r_bits_resp;
  wire[63:0] err_slave_io_r_bits_data;
  wire err_slave_io_r_bits_last;
  wire[4:0] err_slave_io_r_bits_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R29 = {1{$random}};
    R40 = {1{$random}};
    R51 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = r_invalid & io_master_ar_valid;
  assign r_invalid = T1 ^ 1'h1;
  assign T1 = ar_route != 3'h0;
  assign ar_route = T2;
  assign T2 = {T10, T3};
  assign T3 = {T7, T4};
  assign T4 = T6 & T5;
  assign T5 = io_master_ar_bits_addr < 32'h40000000;
  assign T6 = 32'h0 <= io_master_ar_bits_addr;
  assign T7 = T9 & T8;
  assign T8 = io_master_ar_bits_addr < 32'h80000000;
  assign T9 = 32'h40000000 <= io_master_ar_bits_addr;
  assign T10 = T12 & T11;
  assign T11 = T82 < 33'h100000000;
  assign T82 = {1'h0, io_master_ar_bits_addr};
  assign T12 = 32'h80000000 <= io_master_ar_bits_addr;
  assign T13 = w_invalid & io_master_aw_valid;
  assign w_invalid = T14 ^ 1'h1;
  assign T14 = aw_route != 3'h0;
  assign aw_route = T15;
  assign T15 = {T23, T16};
  assign T16 = {T20, T17};
  assign T17 = T19 & T18;
  assign T18 = io_master_aw_bits_addr < 32'h40000000;
  assign T19 = 32'h0 <= io_master_aw_bits_addr;
  assign T20 = T22 & T21;
  assign T21 = io_master_aw_bits_addr < 32'h80000000;
  assign T22 = 32'h40000000 <= io_master_aw_bits_addr;
  assign T23 = T25 & T24;
  assign T24 = T83 < 33'h100000000;
  assign T83 = {1'h0, io_master_aw_bits_addr};
  assign T25 = 32'h80000000 <= io_master_aw_bits_addr;
  assign io_slave_0_r_ready = r_arb_io_in_0_ready;
  assign io_slave_0_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_0_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_0_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_0_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_0_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_0_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_0_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_0_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_0_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_0_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_0_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_0_ar_valid = T26;
  assign T26 = io_master_ar_valid & T27;
  assign T27 = ar_route[1'h0:1'h0];
  assign io_slave_0_b_ready = b_arb_io_in_0_ready;
  assign io_slave_0_w_bits_user = io_master_w_bits_user;
  assign io_slave_0_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_0_w_bits_last = io_master_w_bits_last;
  assign io_slave_0_w_bits_data = io_master_w_bits_data;
  assign io_slave_0_w_valid = T28;
  assign T28 = io_master_w_valid & R29;
  assign T84 = reset ? 1'h0 : T30;
  assign T30 = T33 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : R29;
  assign T32 = io_slave_0_aw_ready & io_slave_0_aw_valid;
  assign T33 = T34 & io_slave_0_w_bits_last;
  assign T34 = io_slave_0_w_ready & io_slave_0_w_valid;
  assign io_slave_0_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_0_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_0_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_0_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_0_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_0_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_0_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_0_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_0_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_0_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_0_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_0_aw_valid = T35;
  assign T35 = io_master_aw_valid & T36;
  assign T36 = aw_route[1'h0:1'h0];
  assign io_slave_1_r_ready = r_arb_io_in_1_ready;
  assign io_slave_1_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_1_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_1_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_1_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_1_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_1_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_1_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_1_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_1_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_1_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_1_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_1_ar_valid = T37;
  assign T37 = io_master_ar_valid & T38;
  assign T38 = ar_route[1'h1:1'h1];
  assign io_slave_1_b_ready = b_arb_io_in_1_ready;
  assign io_slave_1_w_bits_user = io_master_w_bits_user;
  assign io_slave_1_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_1_w_bits_last = io_master_w_bits_last;
  assign io_slave_1_w_bits_data = io_master_w_bits_data;
  assign io_slave_1_w_valid = T39;
  assign T39 = io_master_w_valid & R40;
  assign T85 = reset ? 1'h0 : T41;
  assign T41 = T44 ? 1'h0 : T42;
  assign T42 = T43 ? 1'h1 : R40;
  assign T43 = io_slave_1_aw_ready & io_slave_1_aw_valid;
  assign T44 = T45 & io_slave_1_w_bits_last;
  assign T45 = io_slave_1_w_ready & io_slave_1_w_valid;
  assign io_slave_1_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_1_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_1_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_1_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_1_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_1_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_1_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_1_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_1_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_1_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_1_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_1_aw_valid = T46;
  assign T46 = io_master_aw_valid & T47;
  assign T47 = aw_route[1'h1:1'h1];
  assign io_slave_2_r_ready = r_arb_io_in_2_ready;
  assign io_slave_2_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_2_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_2_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_2_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_2_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_2_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_2_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_2_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_2_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_2_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_2_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_2_ar_valid = T48;
  assign T48 = io_master_ar_valid & T49;
  assign T49 = ar_route[2'h2:2'h2];
  assign io_slave_2_b_ready = b_arb_io_in_2_ready;
  assign io_slave_2_w_bits_user = io_master_w_bits_user;
  assign io_slave_2_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_2_w_bits_last = io_master_w_bits_last;
  assign io_slave_2_w_bits_data = io_master_w_bits_data;
  assign io_slave_2_w_valid = T50;
  assign T50 = io_master_w_valid & R51;
  assign T86 = reset ? 1'h0 : T52;
  assign T52 = T55 ? 1'h0 : T53;
  assign T53 = T54 ? 1'h1 : R51;
  assign T54 = io_slave_2_aw_ready & io_slave_2_aw_valid;
  assign T55 = T56 & io_slave_2_w_bits_last;
  assign T56 = io_slave_2_w_ready & io_slave_2_w_valid;
  assign io_slave_2_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_2_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_2_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_2_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_2_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_2_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_2_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_2_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_2_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_2_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_2_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_2_aw_valid = T57;
  assign T57 = io_master_aw_valid & T58;
  assign T58 = aw_route[2'h2:2'h2];
  assign io_master_r_bits_user = r_arb_io_out_bits_user;
  assign io_master_r_bits_id = r_arb_io_out_bits_id;
  assign io_master_r_bits_last = r_arb_io_out_bits_last;
  assign io_master_r_bits_data = r_arb_io_out_bits_data;
  assign io_master_r_bits_resp = r_arb_io_out_bits_resp;
  assign io_master_r_valid = r_arb_io_out_valid;
  assign io_master_ar_ready = T59;
  assign T59 = ar_ready | T60;
  assign T60 = r_invalid & err_slave_io_ar_ready;
  assign ar_ready = T63 | T61;
  assign T61 = io_slave_2_ar_ready & T62;
  assign T62 = ar_route[2'h2:2'h2];
  assign T63 = T66 | T64;
  assign T64 = io_slave_1_ar_ready & T65;
  assign T65 = ar_route[1'h1:1'h1];
  assign T66 = io_slave_0_ar_ready & T67;
  assign T67 = ar_route[1'h0:1'h0];
  assign io_master_b_bits_user = b_arb_io_out_bits_user;
  assign io_master_b_bits_id = b_arb_io_out_bits_id;
  assign io_master_b_bits_resp = b_arb_io_out_bits_resp;
  assign io_master_b_valid = b_arb_io_out_valid;
  assign io_master_w_ready = T68;
  assign T68 = w_ready | err_slave_io_w_ready;
  assign w_ready = T70 | T69;
  assign T69 = io_slave_2_w_ready & R51;
  assign T70 = T72 | T71;
  assign T71 = io_slave_1_w_ready & R40;
  assign T72 = io_slave_0_w_ready & R29;
  assign io_master_aw_ready = T73;
  assign T73 = aw_ready | T74;
  assign T74 = w_invalid & err_slave_io_aw_ready;
  assign aw_ready = T77 | T75;
  assign T75 = io_slave_2_aw_ready & T76;
  assign T76 = aw_route[2'h2:2'h2];
  assign T77 = T80 | T78;
  assign T78 = io_slave_1_aw_ready & T79;
  assign T79 = aw_route[1'h1:1'h1];
  assign T80 = io_slave_0_aw_ready & T81;
  assign T81 = aw_route[1'h0:1'h0];
  NastiErrorSlave err_slave(.clk(clk), .reset(reset),
       .io_aw_ready( err_slave_io_aw_ready ),
       .io_aw_valid( T13 ),
       .io_aw_bits_addr( io_master_aw_bits_addr ),
       .io_aw_bits_len( io_master_aw_bits_len ),
       .io_aw_bits_size( io_master_aw_bits_size ),
       .io_aw_bits_burst( io_master_aw_bits_burst ),
       .io_aw_bits_lock( io_master_aw_bits_lock ),
       .io_aw_bits_cache( io_master_aw_bits_cache ),
       .io_aw_bits_prot( io_master_aw_bits_prot ),
       .io_aw_bits_qos( io_master_aw_bits_qos ),
       .io_aw_bits_region( io_master_aw_bits_region ),
       .io_aw_bits_id( io_master_aw_bits_id ),
       .io_aw_bits_user( io_master_aw_bits_user ),
       .io_w_ready( err_slave_io_w_ready ),
       .io_w_valid( io_master_w_valid ),
       .io_w_bits_data( io_master_w_bits_data ),
       .io_w_bits_last( io_master_w_bits_last ),
       .io_w_bits_strb( io_master_w_bits_strb ),
       .io_w_bits_user( io_master_w_bits_user ),
       .io_b_ready( b_arb_io_in_3_ready ),
       .io_b_valid( err_slave_io_b_valid ),
       .io_b_bits_resp( err_slave_io_b_bits_resp ),
       .io_b_bits_id( err_slave_io_b_bits_id ),
       //.io_b_bits_user(  )
       .io_ar_ready( err_slave_io_ar_ready ),
       .io_ar_valid( T0 ),
       .io_ar_bits_addr( io_master_ar_bits_addr ),
       .io_ar_bits_len( io_master_ar_bits_len ),
       .io_ar_bits_size( io_master_ar_bits_size ),
       .io_ar_bits_burst( io_master_ar_bits_burst ),
       .io_ar_bits_lock( io_master_ar_bits_lock ),
       .io_ar_bits_cache( io_master_ar_bits_cache ),
       .io_ar_bits_prot( io_master_ar_bits_prot ),
       .io_ar_bits_qos( io_master_ar_bits_qos ),
       .io_ar_bits_region( io_master_ar_bits_region ),
       .io_ar_bits_id( io_master_ar_bits_id ),
       .io_ar_bits_user( io_master_ar_bits_user ),
       .io_r_ready( r_arb_io_in_3_ready ),
       .io_r_valid( err_slave_io_r_valid ),
       .io_r_bits_resp( err_slave_io_r_bits_resp ),
       .io_r_bits_data( err_slave_io_r_bits_data ),
       .io_r_bits_last( err_slave_io_r_bits_last ),
       .io_r_bits_id( err_slave_io_r_bits_id )
       //.io_r_bits_user(  )
  );
  RRArbiter_4 b_arb(.clk(clk), .reset(reset),
       .io_in_3_ready( b_arb_io_in_3_ready ),
       .io_in_3_valid( err_slave_io_b_valid ),
       .io_in_3_bits_resp( err_slave_io_b_bits_resp ),
       .io_in_3_bits_id( err_slave_io_b_bits_id ),
       //.io_in_3_bits_user(  )
       .io_in_2_ready( b_arb_io_in_2_ready ),
       .io_in_2_valid( io_slave_2_b_valid ),
       .io_in_2_bits_resp( io_slave_2_b_bits_resp ),
       .io_in_2_bits_id( io_slave_2_b_bits_id ),
       .io_in_2_bits_user( io_slave_2_b_bits_user ),
       .io_in_1_ready( b_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_b_valid ),
       .io_in_1_bits_resp( io_slave_1_b_bits_resp ),
       .io_in_1_bits_id( io_slave_1_b_bits_id ),
       .io_in_1_bits_user( io_slave_1_b_bits_user ),
       .io_in_0_ready( b_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_b_valid ),
       .io_in_0_bits_resp( io_slave_0_b_bits_resp ),
       .io_in_0_bits_id( io_slave_0_b_bits_id ),
       .io_in_0_bits_user( io_slave_0_b_bits_user ),
       .io_out_ready( io_master_b_ready ),
       .io_out_valid( b_arb_io_out_valid ),
       .io_out_bits_resp( b_arb_io_out_bits_resp ),
       .io_out_bits_id( b_arb_io_out_bits_id ),
       .io_out_bits_user( b_arb_io_out_bits_user )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign b_arb.io_in_3_bits_user = {1{$random}};
// synthesis translate_on
`endif
  JunctionsPeekingArbiter_0 r_arb(.clk(clk), .reset(reset),
       .io_in_3_ready( r_arb_io_in_3_ready ),
       .io_in_3_valid( err_slave_io_r_valid ),
       .io_in_3_bits_resp( err_slave_io_r_bits_resp ),
       .io_in_3_bits_data( err_slave_io_r_bits_data ),
       .io_in_3_bits_last( err_slave_io_r_bits_last ),
       .io_in_3_bits_id( err_slave_io_r_bits_id ),
       //.io_in_3_bits_user(  )
       .io_in_2_ready( r_arb_io_in_2_ready ),
       .io_in_2_valid( io_slave_2_r_valid ),
       .io_in_2_bits_resp( io_slave_2_r_bits_resp ),
       .io_in_2_bits_data( io_slave_2_r_bits_data ),
       .io_in_2_bits_last( io_slave_2_r_bits_last ),
       .io_in_2_bits_id( io_slave_2_r_bits_id ),
       .io_in_2_bits_user( io_slave_2_r_bits_user ),
       .io_in_1_ready( r_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_r_valid ),
       .io_in_1_bits_resp( io_slave_1_r_bits_resp ),
       .io_in_1_bits_data( io_slave_1_r_bits_data ),
       .io_in_1_bits_last( io_slave_1_r_bits_last ),
       .io_in_1_bits_id( io_slave_1_r_bits_id ),
       .io_in_1_bits_user( io_slave_1_r_bits_user ),
       .io_in_0_ready( r_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_r_valid ),
       .io_in_0_bits_resp( io_slave_0_r_bits_resp ),
       .io_in_0_bits_data( io_slave_0_r_bits_data ),
       .io_in_0_bits_last( io_slave_0_r_bits_last ),
       .io_in_0_bits_id( io_slave_0_r_bits_id ),
       .io_in_0_bits_user( io_slave_0_r_bits_user ),
       .io_out_ready( io_master_r_ready ),
       .io_out_valid( r_arb_io_out_valid ),
       .io_out_bits_resp( r_arb_io_out_bits_resp ),
       .io_out_bits_data( r_arb_io_out_bits_data ),
       .io_out_bits_last( r_arb_io_out_bits_last ),
       .io_out_bits_id( r_arb_io_out_bits_id ),
       .io_out_bits_user( r_arb_io_out_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign r_arb.io_in_3_bits_user = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      R29 <= 1'h0;
    end else if(T33) begin
      R29 <= 1'h0;
    end else if(T32) begin
      R29 <= 1'h1;
    end
    if(reset) begin
      R40 <= 1'h0;
    end else if(T44) begin
      R40 <= 1'h0;
    end else if(T43) begin
      R40 <= 1'h1;
    end
    if(reset) begin
      R51 <= 1'h0;
    end else if(T55) begin
      R51 <= 1'h0;
    end else if(T54) begin
      R51 <= 1'h1;
    end
  end
endmodule

module RRArbiter_5(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [31:0] io_in_1_bits_addr,
    input [7:0] io_in_1_bits_len,
    input [2:0] io_in_1_bits_size,
    input [1:0] io_in_1_bits_burst,
    input  io_in_1_bits_lock,
    input [3:0] io_in_1_bits_cache,
    input [2:0] io_in_1_bits_prot,
    input [3:0] io_in_1_bits_qos,
    input [3:0] io_in_1_bits_region,
    input [4:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [31:0] io_in_0_bits_addr,
    input [7:0] io_in_0_bits_len,
    input [2:0] io_in_0_bits_size,
    input [1:0] io_in_0_bits_burst,
    input  io_in_0_bits_lock,
    input [3:0] io_in_0_bits_cache,
    input [2:0] io_in_0_bits_prot,
    input [3:0] io_in_0_bits_qos,
    input [3:0] io_in_0_bits_region,
    input [4:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits_addr,
    output[7:0] io_out_bits_len,
    output[2:0] io_out_bits_size,
    output[1:0] io_out_bits_burst,
    output io_out_bits_lock,
    output[3:0] io_out_bits_cache,
    output[2:0] io_out_bits_prot,
    output[3:0] io_out_bits_qos,
    output[3:0] io_out_bits_region,
    output[4:0] io_out_bits_id,
    output io_out_bits_user,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T35;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[4:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[2:0] T10;
  wire[3:0] T11;
  wire T12;
  wire[1:0] T13;
  wire[2:0] T14;
  wire[7:0] T15;
  wire[31:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T35 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_user = T5;
  assign T5 = T6 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T6 = chosen;
  assign io_out_bits_id = T7;
  assign T7 = T6 ? io_in_1_bits_id : io_in_0_bits_id;
  assign io_out_bits_region = T8;
  assign T8 = T6 ? io_in_1_bits_region : io_in_0_bits_region;
  assign io_out_bits_qos = T9;
  assign T9 = T6 ? io_in_1_bits_qos : io_in_0_bits_qos;
  assign io_out_bits_prot = T10;
  assign T10 = T6 ? io_in_1_bits_prot : io_in_0_bits_prot;
  assign io_out_bits_cache = T11;
  assign T11 = T6 ? io_in_1_bits_cache : io_in_0_bits_cache;
  assign io_out_bits_lock = T12;
  assign T12 = T6 ? io_in_1_bits_lock : io_in_0_bits_lock;
  assign io_out_bits_burst = T13;
  assign T13 = T6 ? io_in_1_bits_burst : io_in_0_bits_burst;
  assign io_out_bits_size = T14;
  assign T14 = T6 ? io_in_1_bits_size : io_in_0_bits_size;
  assign io_out_bits_len = T15;
  assign T15 = T6 ? io_in_1_bits_len : io_in_0_bits_len;
  assign io_out_bits_addr = T16;
  assign T16 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T17;
  assign T17 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T18;
  assign T18 = T19 & io_out_ready;
  assign T19 = T26 | T20;
  assign T20 = T21 ^ 1'h1;
  assign T21 = T24 | T22;
  assign T22 = io_in_1_valid & T23;
  assign T23 = last_grant < 1'h1;
  assign T24 = io_in_0_valid & T25;
  assign T25 = last_grant < 1'h0;
  assign T26 = last_grant < 1'h0;
  assign io_in_1_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T32 | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 | io_in_0_valid;
  assign T31 = T24 | T22;
  assign T32 = T34 & T33;
  assign T33 = last_grant < 1'h1;
  assign T34 = T24 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module NastiArbiter(input clk, input reset,
    output io_master_1_aw_ready,
    input  io_master_1_aw_valid,
    input [31:0] io_master_1_aw_bits_addr,
    input [7:0] io_master_1_aw_bits_len,
    input [2:0] io_master_1_aw_bits_size,
    input [1:0] io_master_1_aw_bits_burst,
    input  io_master_1_aw_bits_lock,
    input [3:0] io_master_1_aw_bits_cache,
    input [2:0] io_master_1_aw_bits_prot,
    input [3:0] io_master_1_aw_bits_qos,
    input [3:0] io_master_1_aw_bits_region,
    input [4:0] io_master_1_aw_bits_id,
    input  io_master_1_aw_bits_user,
    output io_master_1_w_ready,
    input  io_master_1_w_valid,
    input [63:0] io_master_1_w_bits_data,
    input  io_master_1_w_bits_last,
    input [7:0] io_master_1_w_bits_strb,
    input  io_master_1_w_bits_user,
    input  io_master_1_b_ready,
    output io_master_1_b_valid,
    output[1:0] io_master_1_b_bits_resp,
    output[4:0] io_master_1_b_bits_id,
    output io_master_1_b_bits_user,
    output io_master_1_ar_ready,
    input  io_master_1_ar_valid,
    input [31:0] io_master_1_ar_bits_addr,
    input [7:0] io_master_1_ar_bits_len,
    input [2:0] io_master_1_ar_bits_size,
    input [1:0] io_master_1_ar_bits_burst,
    input  io_master_1_ar_bits_lock,
    input [3:0] io_master_1_ar_bits_cache,
    input [2:0] io_master_1_ar_bits_prot,
    input [3:0] io_master_1_ar_bits_qos,
    input [3:0] io_master_1_ar_bits_region,
    input [4:0] io_master_1_ar_bits_id,
    input  io_master_1_ar_bits_user,
    input  io_master_1_r_ready,
    output io_master_1_r_valid,
    output[1:0] io_master_1_r_bits_resp,
    output[63:0] io_master_1_r_bits_data,
    output io_master_1_r_bits_last,
    output[4:0] io_master_1_r_bits_id,
    output io_master_1_r_bits_user,
    output io_master_0_aw_ready,
    input  io_master_0_aw_valid,
    input [31:0] io_master_0_aw_bits_addr,
    input [7:0] io_master_0_aw_bits_len,
    input [2:0] io_master_0_aw_bits_size,
    input [1:0] io_master_0_aw_bits_burst,
    input  io_master_0_aw_bits_lock,
    input [3:0] io_master_0_aw_bits_cache,
    input [2:0] io_master_0_aw_bits_prot,
    input [3:0] io_master_0_aw_bits_qos,
    input [3:0] io_master_0_aw_bits_region,
    input [4:0] io_master_0_aw_bits_id,
    input  io_master_0_aw_bits_user,
    output io_master_0_w_ready,
    input  io_master_0_w_valid,
    input [63:0] io_master_0_w_bits_data,
    input  io_master_0_w_bits_last,
    input [7:0] io_master_0_w_bits_strb,
    input  io_master_0_w_bits_user,
    input  io_master_0_b_ready,
    output io_master_0_b_valid,
    output[1:0] io_master_0_b_bits_resp,
    output[4:0] io_master_0_b_bits_id,
    output io_master_0_b_bits_user,
    output io_master_0_ar_ready,
    input  io_master_0_ar_valid,
    input [31:0] io_master_0_ar_bits_addr,
    input [7:0] io_master_0_ar_bits_len,
    input [2:0] io_master_0_ar_bits_size,
    input [1:0] io_master_0_ar_bits_burst,
    input  io_master_0_ar_bits_lock,
    input [3:0] io_master_0_ar_bits_cache,
    input [2:0] io_master_0_ar_bits_prot,
    input [3:0] io_master_0_ar_bits_qos,
    input [3:0] io_master_0_ar_bits_region,
    input [4:0] io_master_0_ar_bits_id,
    input  io_master_0_ar_bits_user,
    input  io_master_0_r_ready,
    output io_master_0_r_valid,
    output[1:0] io_master_0_r_bits_resp,
    output[63:0] io_master_0_r_bits_data,
    output io_master_0_r_bits_last,
    output[4:0] io_master_0_r_bits_id,
    output io_master_0_r_bits_user,
    input  io_slave_aw_ready,
    output io_slave_aw_valid,
    output[31:0] io_slave_aw_bits_addr,
    output[7:0] io_slave_aw_bits_len,
    output[2:0] io_slave_aw_bits_size,
    output[1:0] io_slave_aw_bits_burst,
    output io_slave_aw_bits_lock,
    output[3:0] io_slave_aw_bits_cache,
    output[2:0] io_slave_aw_bits_prot,
    output[3:0] io_slave_aw_bits_qos,
    output[3:0] io_slave_aw_bits_region,
    output[4:0] io_slave_aw_bits_id,
    output io_slave_aw_bits_user,
    input  io_slave_w_ready,
    output io_slave_w_valid,
    output[63:0] io_slave_w_bits_data,
    output io_slave_w_bits_last,
    output[7:0] io_slave_w_bits_strb,
    output io_slave_w_bits_user,
    output io_slave_b_ready,
    input  io_slave_b_valid,
    input [1:0] io_slave_b_bits_resp,
    input [4:0] io_slave_b_bits_id,
    input  io_slave_b_bits_user,
    input  io_slave_ar_ready,
    output io_slave_ar_valid,
    output[31:0] io_slave_ar_bits_addr,
    output[7:0] io_slave_ar_bits_len,
    output[2:0] io_slave_ar_bits_size,
    output[1:0] io_slave_ar_bits_burst,
    output io_slave_ar_bits_lock,
    output[3:0] io_slave_ar_bits_cache,
    output[2:0] io_slave_ar_bits_prot,
    output[3:0] io_slave_ar_bits_qos,
    output[3:0] io_slave_ar_bits_region,
    output[4:0] io_slave_ar_bits_id,
    output io_slave_ar_bits_user,
    output io_slave_r_ready,
    input  io_slave_r_valid,
    input [1:0] io_slave_r_bits_resp,
    input [63:0] io_slave_r_bits_data,
    input  io_slave_r_bits_last,
    input [4:0] io_slave_r_bits_id,
    input  io_slave_r_bits_user
);

  wire T0;
  reg  R1;
  wire T48;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[4:0] T49;
  wire[5:0] T7;
  wire[4:0] T50;
  wire[5:0] T8;
  wire[4:0] T51;
  wire[5:0] T9;
  wire[4:0] T52;
  wire[5:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg  R19;
  wire T20;
  wire[7:0] T21;
  wire T22;
  wire[63:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[4:0] T53;
  wire[3:0] T28;
  wire T29;
  wire T30;
  wire[4:0] T54;
  wire[3:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[4:0] T55;
  wire[3:0] T38;
  wire T39;
  wire T40;
  wire[4:0] T56;
  wire[3:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire RRArbiter_io_in_1_ready;
  wire RRArbiter_io_in_0_ready;
  wire RRArbiter_io_out_valid;
  wire[31:0] RRArbiter_io_out_bits_addr;
  wire[7:0] RRArbiter_io_out_bits_len;
  wire[2:0] RRArbiter_io_out_bits_size;
  wire[1:0] RRArbiter_io_out_bits_burst;
  wire RRArbiter_io_out_bits_lock;
  wire[3:0] RRArbiter_io_out_bits_cache;
  wire[2:0] RRArbiter_io_out_bits_prot;
  wire[3:0] RRArbiter_io_out_bits_qos;
  wire[3:0] RRArbiter_io_out_bits_region;
  wire[4:0] RRArbiter_io_out_bits_id;
  wire RRArbiter_io_out_bits_user;
  wire RRArbiter_1_io_in_1_ready;
  wire RRArbiter_1_io_in_0_ready;
  wire RRArbiter_1_io_out_valid;
  wire[31:0] RRArbiter_1_io_out_bits_addr;
  wire[7:0] RRArbiter_1_io_out_bits_len;
  wire[2:0] RRArbiter_1_io_out_bits_size;
  wire[1:0] RRArbiter_1_io_out_bits_burst;
  wire RRArbiter_1_io_out_bits_lock;
  wire[3:0] RRArbiter_1_io_out_bits_cache;
  wire[2:0] RRArbiter_1_io_out_bits_prot;
  wire[3:0] RRArbiter_1_io_out_bits_qos;
  wire[3:0] RRArbiter_1_io_out_bits_region;
  wire[4:0] RRArbiter_1_io_out_bits_id;
  wire RRArbiter_1_io_out_bits_user;
  wire RRArbiter_1_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R19 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_slave_aw_ready & R1;
  assign T48 = reset ? 1'h1 : T2;
  assign T2 = T5 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : R1;
  assign T4 = T0 & RRArbiter_1_io_out_valid;
  assign T5 = T6 & io_slave_w_bits_last;
  assign T6 = io_slave_w_ready & io_slave_w_valid;
  assign T49 = T7[3'h4:1'h0];
  assign T7 = {io_master_0_aw_bits_id, 1'h0};
  assign T50 = T8[3'h4:1'h0];
  assign T8 = {io_master_1_aw_bits_id, 1'h1};
  assign T51 = T9[3'h4:1'h0];
  assign T9 = {io_master_0_ar_bits_id, 1'h0};
  assign T52 = T10[3'h4:1'h0];
  assign T10 = {io_master_1_ar_bits_id, 1'h1};
  assign io_slave_r_ready = T11;
  assign T11 = T12 ? io_master_1_r_ready : io_master_0_r_ready;
  assign T12 = T13;
  assign T13 = io_slave_r_bits_id[1'h0:1'h0];
  assign io_slave_ar_bits_user = RRArbiter_io_out_bits_user;
  assign io_slave_ar_bits_id = RRArbiter_io_out_bits_id;
  assign io_slave_ar_bits_region = RRArbiter_io_out_bits_region;
  assign io_slave_ar_bits_qos = RRArbiter_io_out_bits_qos;
  assign io_slave_ar_bits_prot = RRArbiter_io_out_bits_prot;
  assign io_slave_ar_bits_cache = RRArbiter_io_out_bits_cache;
  assign io_slave_ar_bits_lock = RRArbiter_io_out_bits_lock;
  assign io_slave_ar_bits_burst = RRArbiter_io_out_bits_burst;
  assign io_slave_ar_bits_size = RRArbiter_io_out_bits_size;
  assign io_slave_ar_bits_len = RRArbiter_io_out_bits_len;
  assign io_slave_ar_bits_addr = RRArbiter_io_out_bits_addr;
  assign io_slave_ar_valid = RRArbiter_io_out_valid;
  assign io_slave_b_ready = T14;
  assign T14 = T15 ? io_master_1_b_ready : io_master_0_b_ready;
  assign T15 = T16;
  assign T16 = io_slave_b_bits_id[1'h0:1'h0];
  assign io_slave_w_bits_user = T17;
  assign T17 = T18 ? io_master_1_w_bits_user : io_master_0_w_bits_user;
  assign T18 = R19;
  assign T20 = T4 ? RRArbiter_1_io_chosen : R19;
  assign io_slave_w_bits_strb = T21;
  assign T21 = T18 ? io_master_1_w_bits_strb : io_master_0_w_bits_strb;
  assign io_slave_w_bits_last = T22;
  assign T22 = T18 ? io_master_1_w_bits_last : io_master_0_w_bits_last;
  assign io_slave_w_bits_data = T23;
  assign T23 = T18 ? io_master_1_w_bits_data : io_master_0_w_bits_data;
  assign io_slave_w_valid = T24;
  assign T24 = T26 & T25;
  assign T25 = R1 ^ 1'h1;
  assign T26 = T18 ? io_master_1_w_valid : io_master_0_w_valid;
  assign io_slave_aw_bits_user = RRArbiter_1_io_out_bits_user;
  assign io_slave_aw_bits_id = RRArbiter_1_io_out_bits_id;
  assign io_slave_aw_bits_region = RRArbiter_1_io_out_bits_region;
  assign io_slave_aw_bits_qos = RRArbiter_1_io_out_bits_qos;
  assign io_slave_aw_bits_prot = RRArbiter_1_io_out_bits_prot;
  assign io_slave_aw_bits_cache = RRArbiter_1_io_out_bits_cache;
  assign io_slave_aw_bits_lock = RRArbiter_1_io_out_bits_lock;
  assign io_slave_aw_bits_burst = RRArbiter_1_io_out_bits_burst;
  assign io_slave_aw_bits_size = RRArbiter_1_io_out_bits_size;
  assign io_slave_aw_bits_len = RRArbiter_1_io_out_bits_len;
  assign io_slave_aw_bits_addr = RRArbiter_1_io_out_bits_addr;
  assign io_slave_aw_valid = T27;
  assign T27 = RRArbiter_1_io_out_valid & R1;
  assign io_master_0_r_bits_user = io_slave_r_bits_user;
  assign io_master_0_r_bits_id = T53;
  assign T53 = {1'h0, T28};
  assign T28 = io_slave_r_bits_id >> 1'h1;
  assign io_master_0_r_bits_last = io_slave_r_bits_last;
  assign io_master_0_r_bits_data = io_slave_r_bits_data;
  assign io_master_0_r_bits_resp = io_slave_r_bits_resp;
  assign io_master_0_r_valid = T29;
  assign T29 = io_slave_r_valid & T30;
  assign T30 = T13 == 1'h0;
  assign io_master_0_ar_ready = RRArbiter_io_in_0_ready;
  assign io_master_0_b_bits_user = io_slave_b_bits_user;
  assign io_master_0_b_bits_id = T54;
  assign T54 = {1'h0, T31};
  assign T31 = io_slave_b_bits_id >> 1'h1;
  assign io_master_0_b_bits_resp = io_slave_b_bits_resp;
  assign io_master_0_b_valid = T32;
  assign T32 = io_slave_b_valid & T33;
  assign T33 = T16 == 1'h0;
  assign io_master_0_w_ready = T34;
  assign T34 = T36 & T35;
  assign T35 = R1 ^ 1'h1;
  assign T36 = io_slave_w_ready & T37;
  assign T37 = R19 == 1'h0;
  assign io_master_0_aw_ready = RRArbiter_1_io_in_0_ready;
  assign io_master_1_r_bits_user = io_slave_r_bits_user;
  assign io_master_1_r_bits_id = T55;
  assign T55 = {1'h0, T38};
  assign T38 = io_slave_r_bits_id >> 1'h1;
  assign io_master_1_r_bits_last = io_slave_r_bits_last;
  assign io_master_1_r_bits_data = io_slave_r_bits_data;
  assign io_master_1_r_bits_resp = io_slave_r_bits_resp;
  assign io_master_1_r_valid = T39;
  assign T39 = io_slave_r_valid & T40;
  assign T40 = T13 == 1'h1;
  assign io_master_1_ar_ready = RRArbiter_io_in_1_ready;
  assign io_master_1_b_bits_user = io_slave_b_bits_user;
  assign io_master_1_b_bits_id = T56;
  assign T56 = {1'h0, T41};
  assign T41 = io_slave_b_bits_id >> 1'h1;
  assign io_master_1_b_bits_resp = io_slave_b_bits_resp;
  assign io_master_1_b_valid = T42;
  assign T42 = io_slave_b_valid & T43;
  assign T43 = T16 == 1'h1;
  assign io_master_1_w_ready = T44;
  assign T44 = T46 & T45;
  assign T45 = R1 ^ 1'h1;
  assign T46 = io_slave_w_ready & T47;
  assign T47 = R19 == 1'h1;
  assign io_master_1_aw_ready = RRArbiter_1_io_in_1_ready;
  RRArbiter_5 RRArbiter(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_io_in_1_ready ),
       .io_in_1_valid( io_master_1_ar_valid ),
       .io_in_1_bits_addr( io_master_1_ar_bits_addr ),
       .io_in_1_bits_len( io_master_1_ar_bits_len ),
       .io_in_1_bits_size( io_master_1_ar_bits_size ),
       .io_in_1_bits_burst( io_master_1_ar_bits_burst ),
       .io_in_1_bits_lock( io_master_1_ar_bits_lock ),
       .io_in_1_bits_cache( io_master_1_ar_bits_cache ),
       .io_in_1_bits_prot( io_master_1_ar_bits_prot ),
       .io_in_1_bits_qos( io_master_1_ar_bits_qos ),
       .io_in_1_bits_region( io_master_1_ar_bits_region ),
       .io_in_1_bits_id( T52 ),
       .io_in_1_bits_user( io_master_1_ar_bits_user ),
       .io_in_0_ready( RRArbiter_io_in_0_ready ),
       .io_in_0_valid( io_master_0_ar_valid ),
       .io_in_0_bits_addr( io_master_0_ar_bits_addr ),
       .io_in_0_bits_len( io_master_0_ar_bits_len ),
       .io_in_0_bits_size( io_master_0_ar_bits_size ),
       .io_in_0_bits_burst( io_master_0_ar_bits_burst ),
       .io_in_0_bits_lock( io_master_0_ar_bits_lock ),
       .io_in_0_bits_cache( io_master_0_ar_bits_cache ),
       .io_in_0_bits_prot( io_master_0_ar_bits_prot ),
       .io_in_0_bits_qos( io_master_0_ar_bits_qos ),
       .io_in_0_bits_region( io_master_0_ar_bits_region ),
       .io_in_0_bits_id( T51 ),
       .io_in_0_bits_user( io_master_0_ar_bits_user ),
       .io_out_ready( io_slave_ar_ready ),
       .io_out_valid( RRArbiter_io_out_valid ),
       .io_out_bits_addr( RRArbiter_io_out_bits_addr ),
       .io_out_bits_len( RRArbiter_io_out_bits_len ),
       .io_out_bits_size( RRArbiter_io_out_bits_size ),
       .io_out_bits_burst( RRArbiter_io_out_bits_burst ),
       .io_out_bits_lock( RRArbiter_io_out_bits_lock ),
       .io_out_bits_cache( RRArbiter_io_out_bits_cache ),
       .io_out_bits_prot( RRArbiter_io_out_bits_prot ),
       .io_out_bits_qos( RRArbiter_io_out_bits_qos ),
       .io_out_bits_region( RRArbiter_io_out_bits_region ),
       .io_out_bits_id( RRArbiter_io_out_bits_id ),
       .io_out_bits_user( RRArbiter_io_out_bits_user )
       //.io_chosen(  )
  );
  RRArbiter_5 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_master_1_aw_valid ),
       .io_in_1_bits_addr( io_master_1_aw_bits_addr ),
       .io_in_1_bits_len( io_master_1_aw_bits_len ),
       .io_in_1_bits_size( io_master_1_aw_bits_size ),
       .io_in_1_bits_burst( io_master_1_aw_bits_burst ),
       .io_in_1_bits_lock( io_master_1_aw_bits_lock ),
       .io_in_1_bits_cache( io_master_1_aw_bits_cache ),
       .io_in_1_bits_prot( io_master_1_aw_bits_prot ),
       .io_in_1_bits_qos( io_master_1_aw_bits_qos ),
       .io_in_1_bits_region( io_master_1_aw_bits_region ),
       .io_in_1_bits_id( T50 ),
       .io_in_1_bits_user( io_master_1_aw_bits_user ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_master_0_aw_valid ),
       .io_in_0_bits_addr( io_master_0_aw_bits_addr ),
       .io_in_0_bits_len( io_master_0_aw_bits_len ),
       .io_in_0_bits_size( io_master_0_aw_bits_size ),
       .io_in_0_bits_burst( io_master_0_aw_bits_burst ),
       .io_in_0_bits_lock( io_master_0_aw_bits_lock ),
       .io_in_0_bits_cache( io_master_0_aw_bits_cache ),
       .io_in_0_bits_prot( io_master_0_aw_bits_prot ),
       .io_in_0_bits_qos( io_master_0_aw_bits_qos ),
       .io_in_0_bits_region( io_master_0_aw_bits_region ),
       .io_in_0_bits_id( T49 ),
       .io_in_0_bits_user( io_master_0_aw_bits_user ),
       .io_out_ready( T0 ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_addr( RRArbiter_1_io_out_bits_addr ),
       .io_out_bits_len( RRArbiter_1_io_out_bits_len ),
       .io_out_bits_size( RRArbiter_1_io_out_bits_size ),
       .io_out_bits_burst( RRArbiter_1_io_out_bits_burst ),
       .io_out_bits_lock( RRArbiter_1_io_out_bits_lock ),
       .io_out_bits_cache( RRArbiter_1_io_out_bits_cache ),
       .io_out_bits_prot( RRArbiter_1_io_out_bits_prot ),
       .io_out_bits_qos( RRArbiter_1_io_out_bits_qos ),
       .io_out_bits_region( RRArbiter_1_io_out_bits_region ),
       .io_out_bits_id( RRArbiter_1_io_out_bits_id ),
       .io_out_bits_user( RRArbiter_1_io_out_bits_user ),
       .io_chosen( RRArbiter_1_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h1;
    end else if(T5) begin
      R1 <= 1'h1;
    end else if(T4) begin
      R1 <= 1'h0;
    end
    if(T4) begin
      R19 <= RRArbiter_1_io_chosen;
    end
  end
endmodule

module NastiCrossbar_0(input clk, input reset,
    output io_masters_1_aw_ready,
    input  io_masters_1_aw_valid,
    input [31:0] io_masters_1_aw_bits_addr,
    input [7:0] io_masters_1_aw_bits_len,
    input [2:0] io_masters_1_aw_bits_size,
    input [1:0] io_masters_1_aw_bits_burst,
    input  io_masters_1_aw_bits_lock,
    input [3:0] io_masters_1_aw_bits_cache,
    input [2:0] io_masters_1_aw_bits_prot,
    input [3:0] io_masters_1_aw_bits_qos,
    input [3:0] io_masters_1_aw_bits_region,
    input [4:0] io_masters_1_aw_bits_id,
    input  io_masters_1_aw_bits_user,
    output io_masters_1_w_ready,
    input  io_masters_1_w_valid,
    input [63:0] io_masters_1_w_bits_data,
    input  io_masters_1_w_bits_last,
    input [7:0] io_masters_1_w_bits_strb,
    input  io_masters_1_w_bits_user,
    input  io_masters_1_b_ready,
    output io_masters_1_b_valid,
    output[1:0] io_masters_1_b_bits_resp,
    output[4:0] io_masters_1_b_bits_id,
    output io_masters_1_b_bits_user,
    output io_masters_1_ar_ready,
    input  io_masters_1_ar_valid,
    input [31:0] io_masters_1_ar_bits_addr,
    input [7:0] io_masters_1_ar_bits_len,
    input [2:0] io_masters_1_ar_bits_size,
    input [1:0] io_masters_1_ar_bits_burst,
    input  io_masters_1_ar_bits_lock,
    input [3:0] io_masters_1_ar_bits_cache,
    input [2:0] io_masters_1_ar_bits_prot,
    input [3:0] io_masters_1_ar_bits_qos,
    input [3:0] io_masters_1_ar_bits_region,
    input [4:0] io_masters_1_ar_bits_id,
    input  io_masters_1_ar_bits_user,
    input  io_masters_1_r_ready,
    output io_masters_1_r_valid,
    output[1:0] io_masters_1_r_bits_resp,
    output[63:0] io_masters_1_r_bits_data,
    output io_masters_1_r_bits_last,
    output[4:0] io_masters_1_r_bits_id,
    output io_masters_1_r_bits_user,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [4:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[4:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [4:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[4:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_2_aw_ready,
    output io_slaves_2_aw_valid,
    output[31:0] io_slaves_2_aw_bits_addr,
    output[7:0] io_slaves_2_aw_bits_len,
    output[2:0] io_slaves_2_aw_bits_size,
    output[1:0] io_slaves_2_aw_bits_burst,
    output io_slaves_2_aw_bits_lock,
    output[3:0] io_slaves_2_aw_bits_cache,
    output[2:0] io_slaves_2_aw_bits_prot,
    output[3:0] io_slaves_2_aw_bits_qos,
    output[3:0] io_slaves_2_aw_bits_region,
    output[4:0] io_slaves_2_aw_bits_id,
    output io_slaves_2_aw_bits_user,
    input  io_slaves_2_w_ready,
    output io_slaves_2_w_valid,
    output[63:0] io_slaves_2_w_bits_data,
    output io_slaves_2_w_bits_last,
    output[7:0] io_slaves_2_w_bits_strb,
    output io_slaves_2_w_bits_user,
    output io_slaves_2_b_ready,
    input  io_slaves_2_b_valid,
    input [1:0] io_slaves_2_b_bits_resp,
    input [4:0] io_slaves_2_b_bits_id,
    input  io_slaves_2_b_bits_user,
    input  io_slaves_2_ar_ready,
    output io_slaves_2_ar_valid,
    output[31:0] io_slaves_2_ar_bits_addr,
    output[7:0] io_slaves_2_ar_bits_len,
    output[2:0] io_slaves_2_ar_bits_size,
    output[1:0] io_slaves_2_ar_bits_burst,
    output io_slaves_2_ar_bits_lock,
    output[3:0] io_slaves_2_ar_bits_cache,
    output[2:0] io_slaves_2_ar_bits_prot,
    output[3:0] io_slaves_2_ar_bits_qos,
    output[3:0] io_slaves_2_ar_bits_region,
    output[4:0] io_slaves_2_ar_bits_id,
    output io_slaves_2_ar_bits_user,
    output io_slaves_2_r_ready,
    input  io_slaves_2_r_valid,
    input [1:0] io_slaves_2_r_bits_resp,
    input [63:0] io_slaves_2_r_bits_data,
    input  io_slaves_2_r_bits_last,
    input [4:0] io_slaves_2_r_bits_id,
    input  io_slaves_2_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[4:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [4:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[4:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [4:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[4:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [4:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[4:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [4:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire NastiArbiter_io_master_1_aw_ready;
  wire NastiArbiter_io_master_1_w_ready;
  wire NastiArbiter_io_master_1_b_valid;
  wire[1:0] NastiArbiter_io_master_1_b_bits_resp;
  wire[4:0] NastiArbiter_io_master_1_b_bits_id;
  wire NastiArbiter_io_master_1_b_bits_user;
  wire NastiArbiter_io_master_1_ar_ready;
  wire NastiArbiter_io_master_1_r_valid;
  wire[1:0] NastiArbiter_io_master_1_r_bits_resp;
  wire[63:0] NastiArbiter_io_master_1_r_bits_data;
  wire NastiArbiter_io_master_1_r_bits_last;
  wire[4:0] NastiArbiter_io_master_1_r_bits_id;
  wire NastiArbiter_io_master_1_r_bits_user;
  wire NastiArbiter_io_master_0_aw_ready;
  wire NastiArbiter_io_master_0_w_ready;
  wire NastiArbiter_io_master_0_b_valid;
  wire[1:0] NastiArbiter_io_master_0_b_bits_resp;
  wire[4:0] NastiArbiter_io_master_0_b_bits_id;
  wire NastiArbiter_io_master_0_b_bits_user;
  wire NastiArbiter_io_master_0_ar_ready;
  wire NastiArbiter_io_master_0_r_valid;
  wire[1:0] NastiArbiter_io_master_0_r_bits_resp;
  wire[63:0] NastiArbiter_io_master_0_r_bits_data;
  wire NastiArbiter_io_master_0_r_bits_last;
  wire[4:0] NastiArbiter_io_master_0_r_bits_id;
  wire NastiArbiter_io_master_0_r_bits_user;
  wire NastiArbiter_io_slave_aw_valid;
  wire[31:0] NastiArbiter_io_slave_aw_bits_addr;
  wire[7:0] NastiArbiter_io_slave_aw_bits_len;
  wire[2:0] NastiArbiter_io_slave_aw_bits_size;
  wire[1:0] NastiArbiter_io_slave_aw_bits_burst;
  wire NastiArbiter_io_slave_aw_bits_lock;
  wire[3:0] NastiArbiter_io_slave_aw_bits_cache;
  wire[2:0] NastiArbiter_io_slave_aw_bits_prot;
  wire[3:0] NastiArbiter_io_slave_aw_bits_qos;
  wire[3:0] NastiArbiter_io_slave_aw_bits_region;
  wire[4:0] NastiArbiter_io_slave_aw_bits_id;
  wire NastiArbiter_io_slave_aw_bits_user;
  wire NastiArbiter_io_slave_w_valid;
  wire[63:0] NastiArbiter_io_slave_w_bits_data;
  wire NastiArbiter_io_slave_w_bits_last;
  wire[7:0] NastiArbiter_io_slave_w_bits_strb;
  wire NastiArbiter_io_slave_w_bits_user;
  wire NastiArbiter_io_slave_b_ready;
  wire NastiArbiter_io_slave_ar_valid;
  wire[31:0] NastiArbiter_io_slave_ar_bits_addr;
  wire[7:0] NastiArbiter_io_slave_ar_bits_len;
  wire[2:0] NastiArbiter_io_slave_ar_bits_size;
  wire[1:0] NastiArbiter_io_slave_ar_bits_burst;
  wire NastiArbiter_io_slave_ar_bits_lock;
  wire[3:0] NastiArbiter_io_slave_ar_bits_cache;
  wire[2:0] NastiArbiter_io_slave_ar_bits_prot;
  wire[3:0] NastiArbiter_io_slave_ar_bits_qos;
  wire[3:0] NastiArbiter_io_slave_ar_bits_region;
  wire[4:0] NastiArbiter_io_slave_ar_bits_id;
  wire NastiArbiter_io_slave_ar_bits_user;
  wire NastiArbiter_io_slave_r_ready;
  wire NastiArbiter_1_io_master_1_aw_ready;
  wire NastiArbiter_1_io_master_1_w_ready;
  wire NastiArbiter_1_io_master_1_b_valid;
  wire[1:0] NastiArbiter_1_io_master_1_b_bits_resp;
  wire[4:0] NastiArbiter_1_io_master_1_b_bits_id;
  wire NastiArbiter_1_io_master_1_b_bits_user;
  wire NastiArbiter_1_io_master_1_ar_ready;
  wire NastiArbiter_1_io_master_1_r_valid;
  wire[1:0] NastiArbiter_1_io_master_1_r_bits_resp;
  wire[63:0] NastiArbiter_1_io_master_1_r_bits_data;
  wire NastiArbiter_1_io_master_1_r_bits_last;
  wire[4:0] NastiArbiter_1_io_master_1_r_bits_id;
  wire NastiArbiter_1_io_master_1_r_bits_user;
  wire NastiArbiter_1_io_master_0_aw_ready;
  wire NastiArbiter_1_io_master_0_w_ready;
  wire NastiArbiter_1_io_master_0_b_valid;
  wire[1:0] NastiArbiter_1_io_master_0_b_bits_resp;
  wire[4:0] NastiArbiter_1_io_master_0_b_bits_id;
  wire NastiArbiter_1_io_master_0_b_bits_user;
  wire NastiArbiter_1_io_master_0_ar_ready;
  wire NastiArbiter_1_io_master_0_r_valid;
  wire[1:0] NastiArbiter_1_io_master_0_r_bits_resp;
  wire[63:0] NastiArbiter_1_io_master_0_r_bits_data;
  wire NastiArbiter_1_io_master_0_r_bits_last;
  wire[4:0] NastiArbiter_1_io_master_0_r_bits_id;
  wire NastiArbiter_1_io_master_0_r_bits_user;
  wire NastiArbiter_1_io_slave_aw_valid;
  wire[31:0] NastiArbiter_1_io_slave_aw_bits_addr;
  wire[7:0] NastiArbiter_1_io_slave_aw_bits_len;
  wire[2:0] NastiArbiter_1_io_slave_aw_bits_size;
  wire[1:0] NastiArbiter_1_io_slave_aw_bits_burst;
  wire NastiArbiter_1_io_slave_aw_bits_lock;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_cache;
  wire[2:0] NastiArbiter_1_io_slave_aw_bits_prot;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_qos;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_region;
  wire[4:0] NastiArbiter_1_io_slave_aw_bits_id;
  wire NastiArbiter_1_io_slave_aw_bits_user;
  wire NastiArbiter_1_io_slave_w_valid;
  wire[63:0] NastiArbiter_1_io_slave_w_bits_data;
  wire NastiArbiter_1_io_slave_w_bits_last;
  wire[7:0] NastiArbiter_1_io_slave_w_bits_strb;
  wire NastiArbiter_1_io_slave_w_bits_user;
  wire NastiArbiter_1_io_slave_b_ready;
  wire NastiArbiter_1_io_slave_ar_valid;
  wire[31:0] NastiArbiter_1_io_slave_ar_bits_addr;
  wire[7:0] NastiArbiter_1_io_slave_ar_bits_len;
  wire[2:0] NastiArbiter_1_io_slave_ar_bits_size;
  wire[1:0] NastiArbiter_1_io_slave_ar_bits_burst;
  wire NastiArbiter_1_io_slave_ar_bits_lock;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_cache;
  wire[2:0] NastiArbiter_1_io_slave_ar_bits_prot;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_qos;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_region;
  wire[4:0] NastiArbiter_1_io_slave_ar_bits_id;
  wire NastiArbiter_1_io_slave_ar_bits_user;
  wire NastiArbiter_1_io_slave_r_ready;
  wire NastiArbiter_2_io_master_1_aw_ready;
  wire NastiArbiter_2_io_master_1_w_ready;
  wire NastiArbiter_2_io_master_1_b_valid;
  wire[1:0] NastiArbiter_2_io_master_1_b_bits_resp;
  wire[4:0] NastiArbiter_2_io_master_1_b_bits_id;
  wire NastiArbiter_2_io_master_1_b_bits_user;
  wire NastiArbiter_2_io_master_1_ar_ready;
  wire NastiArbiter_2_io_master_1_r_valid;
  wire[1:0] NastiArbiter_2_io_master_1_r_bits_resp;
  wire[63:0] NastiArbiter_2_io_master_1_r_bits_data;
  wire NastiArbiter_2_io_master_1_r_bits_last;
  wire[4:0] NastiArbiter_2_io_master_1_r_bits_id;
  wire NastiArbiter_2_io_master_1_r_bits_user;
  wire NastiArbiter_2_io_master_0_aw_ready;
  wire NastiArbiter_2_io_master_0_w_ready;
  wire NastiArbiter_2_io_master_0_b_valid;
  wire[1:0] NastiArbiter_2_io_master_0_b_bits_resp;
  wire[4:0] NastiArbiter_2_io_master_0_b_bits_id;
  wire NastiArbiter_2_io_master_0_b_bits_user;
  wire NastiArbiter_2_io_master_0_ar_ready;
  wire NastiArbiter_2_io_master_0_r_valid;
  wire[1:0] NastiArbiter_2_io_master_0_r_bits_resp;
  wire[63:0] NastiArbiter_2_io_master_0_r_bits_data;
  wire NastiArbiter_2_io_master_0_r_bits_last;
  wire[4:0] NastiArbiter_2_io_master_0_r_bits_id;
  wire NastiArbiter_2_io_master_0_r_bits_user;
  wire NastiArbiter_2_io_slave_aw_valid;
  wire[31:0] NastiArbiter_2_io_slave_aw_bits_addr;
  wire[7:0] NastiArbiter_2_io_slave_aw_bits_len;
  wire[2:0] NastiArbiter_2_io_slave_aw_bits_size;
  wire[1:0] NastiArbiter_2_io_slave_aw_bits_burst;
  wire NastiArbiter_2_io_slave_aw_bits_lock;
  wire[3:0] NastiArbiter_2_io_slave_aw_bits_cache;
  wire[2:0] NastiArbiter_2_io_slave_aw_bits_prot;
  wire[3:0] NastiArbiter_2_io_slave_aw_bits_qos;
  wire[3:0] NastiArbiter_2_io_slave_aw_bits_region;
  wire[4:0] NastiArbiter_2_io_slave_aw_bits_id;
  wire NastiArbiter_2_io_slave_aw_bits_user;
  wire NastiArbiter_2_io_slave_w_valid;
  wire[63:0] NastiArbiter_2_io_slave_w_bits_data;
  wire NastiArbiter_2_io_slave_w_bits_last;
  wire[7:0] NastiArbiter_2_io_slave_w_bits_strb;
  wire NastiArbiter_2_io_slave_w_bits_user;
  wire NastiArbiter_2_io_slave_b_ready;
  wire NastiArbiter_2_io_slave_ar_valid;
  wire[31:0] NastiArbiter_2_io_slave_ar_bits_addr;
  wire[7:0] NastiArbiter_2_io_slave_ar_bits_len;
  wire[2:0] NastiArbiter_2_io_slave_ar_bits_size;
  wire[1:0] NastiArbiter_2_io_slave_ar_bits_burst;
  wire NastiArbiter_2_io_slave_ar_bits_lock;
  wire[3:0] NastiArbiter_2_io_slave_ar_bits_cache;
  wire[2:0] NastiArbiter_2_io_slave_ar_bits_prot;
  wire[3:0] NastiArbiter_2_io_slave_ar_bits_qos;
  wire[3:0] NastiArbiter_2_io_slave_ar_bits_region;
  wire[4:0] NastiArbiter_2_io_slave_ar_bits_id;
  wire NastiArbiter_2_io_slave_ar_bits_user;
  wire NastiArbiter_2_io_slave_r_ready;
  wire NastiRouter_io_master_aw_ready;
  wire NastiRouter_io_master_w_ready;
  wire NastiRouter_io_master_b_valid;
  wire[1:0] NastiRouter_io_master_b_bits_resp;
  wire[4:0] NastiRouter_io_master_b_bits_id;
  wire NastiRouter_io_master_b_bits_user;
  wire NastiRouter_io_master_ar_ready;
  wire NastiRouter_io_master_r_valid;
  wire[1:0] NastiRouter_io_master_r_bits_resp;
  wire[63:0] NastiRouter_io_master_r_bits_data;
  wire NastiRouter_io_master_r_bits_last;
  wire[4:0] NastiRouter_io_master_r_bits_id;
  wire NastiRouter_io_master_r_bits_user;
  wire NastiRouter_io_slave_2_aw_valid;
  wire[31:0] NastiRouter_io_slave_2_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_2_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_2_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_2_aw_bits_burst;
  wire NastiRouter_io_slave_2_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_2_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_region;
  wire[4:0] NastiRouter_io_slave_2_aw_bits_id;
  wire NastiRouter_io_slave_2_aw_bits_user;
  wire NastiRouter_io_slave_2_w_valid;
  wire[63:0] NastiRouter_io_slave_2_w_bits_data;
  wire NastiRouter_io_slave_2_w_bits_last;
  wire[7:0] NastiRouter_io_slave_2_w_bits_strb;
  wire NastiRouter_io_slave_2_w_bits_user;
  wire NastiRouter_io_slave_2_b_ready;
  wire NastiRouter_io_slave_2_ar_valid;
  wire[31:0] NastiRouter_io_slave_2_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_2_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_2_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_2_ar_bits_burst;
  wire NastiRouter_io_slave_2_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_2_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_region;
  wire[4:0] NastiRouter_io_slave_2_ar_bits_id;
  wire NastiRouter_io_slave_2_ar_bits_user;
  wire NastiRouter_io_slave_2_r_ready;
  wire NastiRouter_io_slave_1_aw_valid;
  wire[31:0] NastiRouter_io_slave_1_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_1_aw_bits_burst;
  wire NastiRouter_io_slave_1_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_region;
  wire[4:0] NastiRouter_io_slave_1_aw_bits_id;
  wire NastiRouter_io_slave_1_aw_bits_user;
  wire NastiRouter_io_slave_1_w_valid;
  wire[63:0] NastiRouter_io_slave_1_w_bits_data;
  wire NastiRouter_io_slave_1_w_bits_last;
  wire[7:0] NastiRouter_io_slave_1_w_bits_strb;
  wire NastiRouter_io_slave_1_w_bits_user;
  wire NastiRouter_io_slave_1_b_ready;
  wire NastiRouter_io_slave_1_ar_valid;
  wire[31:0] NastiRouter_io_slave_1_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_1_ar_bits_burst;
  wire NastiRouter_io_slave_1_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_region;
  wire[4:0] NastiRouter_io_slave_1_ar_bits_id;
  wire NastiRouter_io_slave_1_ar_bits_user;
  wire NastiRouter_io_slave_1_r_ready;
  wire NastiRouter_io_slave_0_aw_valid;
  wire[31:0] NastiRouter_io_slave_0_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_0_aw_bits_burst;
  wire NastiRouter_io_slave_0_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_region;
  wire[4:0] NastiRouter_io_slave_0_aw_bits_id;
  wire NastiRouter_io_slave_0_aw_bits_user;
  wire NastiRouter_io_slave_0_w_valid;
  wire[63:0] NastiRouter_io_slave_0_w_bits_data;
  wire NastiRouter_io_slave_0_w_bits_last;
  wire[7:0] NastiRouter_io_slave_0_w_bits_strb;
  wire NastiRouter_io_slave_0_w_bits_user;
  wire NastiRouter_io_slave_0_b_ready;
  wire NastiRouter_io_slave_0_ar_valid;
  wire[31:0] NastiRouter_io_slave_0_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_0_ar_bits_burst;
  wire NastiRouter_io_slave_0_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_region;
  wire[4:0] NastiRouter_io_slave_0_ar_bits_id;
  wire NastiRouter_io_slave_0_ar_bits_user;
  wire NastiRouter_io_slave_0_r_ready;
  wire NastiRouter_1_io_master_aw_ready;
  wire NastiRouter_1_io_master_w_ready;
  wire NastiRouter_1_io_master_b_valid;
  wire[1:0] NastiRouter_1_io_master_b_bits_resp;
  wire[4:0] NastiRouter_1_io_master_b_bits_id;
  wire NastiRouter_1_io_master_b_bits_user;
  wire NastiRouter_1_io_master_ar_ready;
  wire NastiRouter_1_io_master_r_valid;
  wire[1:0] NastiRouter_1_io_master_r_bits_resp;
  wire[63:0] NastiRouter_1_io_master_r_bits_data;
  wire NastiRouter_1_io_master_r_bits_last;
  wire[4:0] NastiRouter_1_io_master_r_bits_id;
  wire NastiRouter_1_io_master_r_bits_user;
  wire NastiRouter_1_io_slave_2_aw_valid;
  wire[31:0] NastiRouter_1_io_slave_2_aw_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_2_aw_bits_len;
  wire[2:0] NastiRouter_1_io_slave_2_aw_bits_size;
  wire[1:0] NastiRouter_1_io_slave_2_aw_bits_burst;
  wire NastiRouter_1_io_slave_2_aw_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_2_aw_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_2_aw_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_2_aw_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_2_aw_bits_region;
  wire[4:0] NastiRouter_1_io_slave_2_aw_bits_id;
  wire NastiRouter_1_io_slave_2_aw_bits_user;
  wire NastiRouter_1_io_slave_2_w_valid;
  wire[63:0] NastiRouter_1_io_slave_2_w_bits_data;
  wire NastiRouter_1_io_slave_2_w_bits_last;
  wire[7:0] NastiRouter_1_io_slave_2_w_bits_strb;
  wire NastiRouter_1_io_slave_2_w_bits_user;
  wire NastiRouter_1_io_slave_2_b_ready;
  wire NastiRouter_1_io_slave_2_ar_valid;
  wire[31:0] NastiRouter_1_io_slave_2_ar_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_2_ar_bits_len;
  wire[2:0] NastiRouter_1_io_slave_2_ar_bits_size;
  wire[1:0] NastiRouter_1_io_slave_2_ar_bits_burst;
  wire NastiRouter_1_io_slave_2_ar_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_2_ar_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_2_ar_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_2_ar_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_2_ar_bits_region;
  wire[4:0] NastiRouter_1_io_slave_2_ar_bits_id;
  wire NastiRouter_1_io_slave_2_ar_bits_user;
  wire NastiRouter_1_io_slave_2_r_ready;
  wire NastiRouter_1_io_slave_1_aw_valid;
  wire[31:0] NastiRouter_1_io_slave_1_aw_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_1_aw_bits_len;
  wire[2:0] NastiRouter_1_io_slave_1_aw_bits_size;
  wire[1:0] NastiRouter_1_io_slave_1_aw_bits_burst;
  wire NastiRouter_1_io_slave_1_aw_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_1_aw_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_region;
  wire[4:0] NastiRouter_1_io_slave_1_aw_bits_id;
  wire NastiRouter_1_io_slave_1_aw_bits_user;
  wire NastiRouter_1_io_slave_1_w_valid;
  wire[63:0] NastiRouter_1_io_slave_1_w_bits_data;
  wire NastiRouter_1_io_slave_1_w_bits_last;
  wire[7:0] NastiRouter_1_io_slave_1_w_bits_strb;
  wire NastiRouter_1_io_slave_1_w_bits_user;
  wire NastiRouter_1_io_slave_1_b_ready;
  wire NastiRouter_1_io_slave_1_ar_valid;
  wire[31:0] NastiRouter_1_io_slave_1_ar_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_1_ar_bits_len;
  wire[2:0] NastiRouter_1_io_slave_1_ar_bits_size;
  wire[1:0] NastiRouter_1_io_slave_1_ar_bits_burst;
  wire NastiRouter_1_io_slave_1_ar_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_1_ar_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_region;
  wire[4:0] NastiRouter_1_io_slave_1_ar_bits_id;
  wire NastiRouter_1_io_slave_1_ar_bits_user;
  wire NastiRouter_1_io_slave_1_r_ready;
  wire NastiRouter_1_io_slave_0_aw_valid;
  wire[31:0] NastiRouter_1_io_slave_0_aw_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_0_aw_bits_len;
  wire[2:0] NastiRouter_1_io_slave_0_aw_bits_size;
  wire[1:0] NastiRouter_1_io_slave_0_aw_bits_burst;
  wire NastiRouter_1_io_slave_0_aw_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_0_aw_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_region;
  wire[4:0] NastiRouter_1_io_slave_0_aw_bits_id;
  wire NastiRouter_1_io_slave_0_aw_bits_user;
  wire NastiRouter_1_io_slave_0_w_valid;
  wire[63:0] NastiRouter_1_io_slave_0_w_bits_data;
  wire NastiRouter_1_io_slave_0_w_bits_last;
  wire[7:0] NastiRouter_1_io_slave_0_w_bits_strb;
  wire NastiRouter_1_io_slave_0_w_bits_user;
  wire NastiRouter_1_io_slave_0_b_ready;
  wire NastiRouter_1_io_slave_0_ar_valid;
  wire[31:0] NastiRouter_1_io_slave_0_ar_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_0_ar_bits_len;
  wire[2:0] NastiRouter_1_io_slave_0_ar_bits_size;
  wire[1:0] NastiRouter_1_io_slave_0_ar_bits_burst;
  wire NastiRouter_1_io_slave_0_ar_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_0_ar_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_region;
  wire[4:0] NastiRouter_1_io_slave_0_ar_bits_id;
  wire NastiRouter_1_io_slave_0_ar_bits_user;
  wire NastiRouter_1_io_slave_0_r_ready;


  assign io_slaves_0_r_ready = NastiArbiter_io_slave_r_ready;
  assign io_slaves_0_ar_bits_user = NastiArbiter_io_slave_ar_bits_user;
  assign io_slaves_0_ar_bits_id = NastiArbiter_io_slave_ar_bits_id;
  assign io_slaves_0_ar_bits_region = NastiArbiter_io_slave_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = NastiArbiter_io_slave_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = NastiArbiter_io_slave_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = NastiArbiter_io_slave_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = NastiArbiter_io_slave_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = NastiArbiter_io_slave_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = NastiArbiter_io_slave_ar_bits_size;
  assign io_slaves_0_ar_bits_len = NastiArbiter_io_slave_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = NastiArbiter_io_slave_ar_bits_addr;
  assign io_slaves_0_ar_valid = NastiArbiter_io_slave_ar_valid;
  assign io_slaves_0_b_ready = NastiArbiter_io_slave_b_ready;
  assign io_slaves_0_w_bits_user = NastiArbiter_io_slave_w_bits_user;
  assign io_slaves_0_w_bits_strb = NastiArbiter_io_slave_w_bits_strb;
  assign io_slaves_0_w_bits_last = NastiArbiter_io_slave_w_bits_last;
  assign io_slaves_0_w_bits_data = NastiArbiter_io_slave_w_bits_data;
  assign io_slaves_0_w_valid = NastiArbiter_io_slave_w_valid;
  assign io_slaves_0_aw_bits_user = NastiArbiter_io_slave_aw_bits_user;
  assign io_slaves_0_aw_bits_id = NastiArbiter_io_slave_aw_bits_id;
  assign io_slaves_0_aw_bits_region = NastiArbiter_io_slave_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = NastiArbiter_io_slave_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = NastiArbiter_io_slave_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = NastiArbiter_io_slave_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = NastiArbiter_io_slave_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = NastiArbiter_io_slave_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = NastiArbiter_io_slave_aw_bits_size;
  assign io_slaves_0_aw_bits_len = NastiArbiter_io_slave_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = NastiArbiter_io_slave_aw_bits_addr;
  assign io_slaves_0_aw_valid = NastiArbiter_io_slave_aw_valid;
  assign io_slaves_1_r_ready = NastiArbiter_1_io_slave_r_ready;
  assign io_slaves_1_ar_bits_user = NastiArbiter_1_io_slave_ar_bits_user;
  assign io_slaves_1_ar_bits_id = NastiArbiter_1_io_slave_ar_bits_id;
  assign io_slaves_1_ar_bits_region = NastiArbiter_1_io_slave_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = NastiArbiter_1_io_slave_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = NastiArbiter_1_io_slave_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = NastiArbiter_1_io_slave_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = NastiArbiter_1_io_slave_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = NastiArbiter_1_io_slave_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = NastiArbiter_1_io_slave_ar_bits_size;
  assign io_slaves_1_ar_bits_len = NastiArbiter_1_io_slave_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = NastiArbiter_1_io_slave_ar_bits_addr;
  assign io_slaves_1_ar_valid = NastiArbiter_1_io_slave_ar_valid;
  assign io_slaves_1_b_ready = NastiArbiter_1_io_slave_b_ready;
  assign io_slaves_1_w_bits_user = NastiArbiter_1_io_slave_w_bits_user;
  assign io_slaves_1_w_bits_strb = NastiArbiter_1_io_slave_w_bits_strb;
  assign io_slaves_1_w_bits_last = NastiArbiter_1_io_slave_w_bits_last;
  assign io_slaves_1_w_bits_data = NastiArbiter_1_io_slave_w_bits_data;
  assign io_slaves_1_w_valid = NastiArbiter_1_io_slave_w_valid;
  assign io_slaves_1_aw_bits_user = NastiArbiter_1_io_slave_aw_bits_user;
  assign io_slaves_1_aw_bits_id = NastiArbiter_1_io_slave_aw_bits_id;
  assign io_slaves_1_aw_bits_region = NastiArbiter_1_io_slave_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = NastiArbiter_1_io_slave_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = NastiArbiter_1_io_slave_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = NastiArbiter_1_io_slave_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = NastiArbiter_1_io_slave_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = NastiArbiter_1_io_slave_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = NastiArbiter_1_io_slave_aw_bits_size;
  assign io_slaves_1_aw_bits_len = NastiArbiter_1_io_slave_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = NastiArbiter_1_io_slave_aw_bits_addr;
  assign io_slaves_1_aw_valid = NastiArbiter_1_io_slave_aw_valid;
  assign io_slaves_2_r_ready = NastiArbiter_2_io_slave_r_ready;
  assign io_slaves_2_ar_bits_user = NastiArbiter_2_io_slave_ar_bits_user;
  assign io_slaves_2_ar_bits_id = NastiArbiter_2_io_slave_ar_bits_id;
  assign io_slaves_2_ar_bits_region = NastiArbiter_2_io_slave_ar_bits_region;
  assign io_slaves_2_ar_bits_qos = NastiArbiter_2_io_slave_ar_bits_qos;
  assign io_slaves_2_ar_bits_prot = NastiArbiter_2_io_slave_ar_bits_prot;
  assign io_slaves_2_ar_bits_cache = NastiArbiter_2_io_slave_ar_bits_cache;
  assign io_slaves_2_ar_bits_lock = NastiArbiter_2_io_slave_ar_bits_lock;
  assign io_slaves_2_ar_bits_burst = NastiArbiter_2_io_slave_ar_bits_burst;
  assign io_slaves_2_ar_bits_size = NastiArbiter_2_io_slave_ar_bits_size;
  assign io_slaves_2_ar_bits_len = NastiArbiter_2_io_slave_ar_bits_len;
  assign io_slaves_2_ar_bits_addr = NastiArbiter_2_io_slave_ar_bits_addr;
  assign io_slaves_2_ar_valid = NastiArbiter_2_io_slave_ar_valid;
  assign io_slaves_2_b_ready = NastiArbiter_2_io_slave_b_ready;
  assign io_slaves_2_w_bits_user = NastiArbiter_2_io_slave_w_bits_user;
  assign io_slaves_2_w_bits_strb = NastiArbiter_2_io_slave_w_bits_strb;
  assign io_slaves_2_w_bits_last = NastiArbiter_2_io_slave_w_bits_last;
  assign io_slaves_2_w_bits_data = NastiArbiter_2_io_slave_w_bits_data;
  assign io_slaves_2_w_valid = NastiArbiter_2_io_slave_w_valid;
  assign io_slaves_2_aw_bits_user = NastiArbiter_2_io_slave_aw_bits_user;
  assign io_slaves_2_aw_bits_id = NastiArbiter_2_io_slave_aw_bits_id;
  assign io_slaves_2_aw_bits_region = NastiArbiter_2_io_slave_aw_bits_region;
  assign io_slaves_2_aw_bits_qos = NastiArbiter_2_io_slave_aw_bits_qos;
  assign io_slaves_2_aw_bits_prot = NastiArbiter_2_io_slave_aw_bits_prot;
  assign io_slaves_2_aw_bits_cache = NastiArbiter_2_io_slave_aw_bits_cache;
  assign io_slaves_2_aw_bits_lock = NastiArbiter_2_io_slave_aw_bits_lock;
  assign io_slaves_2_aw_bits_burst = NastiArbiter_2_io_slave_aw_bits_burst;
  assign io_slaves_2_aw_bits_size = NastiArbiter_2_io_slave_aw_bits_size;
  assign io_slaves_2_aw_bits_len = NastiArbiter_2_io_slave_aw_bits_len;
  assign io_slaves_2_aw_bits_addr = NastiArbiter_2_io_slave_aw_bits_addr;
  assign io_slaves_2_aw_valid = NastiArbiter_2_io_slave_aw_valid;
  assign io_masters_0_r_bits_user = NastiRouter_io_master_r_bits_user;
  assign io_masters_0_r_bits_id = NastiRouter_io_master_r_bits_id;
  assign io_masters_0_r_bits_last = NastiRouter_io_master_r_bits_last;
  assign io_masters_0_r_bits_data = NastiRouter_io_master_r_bits_data;
  assign io_masters_0_r_bits_resp = NastiRouter_io_master_r_bits_resp;
  assign io_masters_0_r_valid = NastiRouter_io_master_r_valid;
  assign io_masters_0_ar_ready = NastiRouter_io_master_ar_ready;
  assign io_masters_0_b_bits_user = NastiRouter_io_master_b_bits_user;
  assign io_masters_0_b_bits_id = NastiRouter_io_master_b_bits_id;
  assign io_masters_0_b_bits_resp = NastiRouter_io_master_b_bits_resp;
  assign io_masters_0_b_valid = NastiRouter_io_master_b_valid;
  assign io_masters_0_w_ready = NastiRouter_io_master_w_ready;
  assign io_masters_0_aw_ready = NastiRouter_io_master_aw_ready;
  assign io_masters_1_r_bits_user = NastiRouter_1_io_master_r_bits_user;
  assign io_masters_1_r_bits_id = NastiRouter_1_io_master_r_bits_id;
  assign io_masters_1_r_bits_last = NastiRouter_1_io_master_r_bits_last;
  assign io_masters_1_r_bits_data = NastiRouter_1_io_master_r_bits_data;
  assign io_masters_1_r_bits_resp = NastiRouter_1_io_master_r_bits_resp;
  assign io_masters_1_r_valid = NastiRouter_1_io_master_r_valid;
  assign io_masters_1_ar_ready = NastiRouter_1_io_master_ar_ready;
  assign io_masters_1_b_bits_user = NastiRouter_1_io_master_b_bits_user;
  assign io_masters_1_b_bits_id = NastiRouter_1_io_master_b_bits_id;
  assign io_masters_1_b_bits_resp = NastiRouter_1_io_master_b_bits_resp;
  assign io_masters_1_b_valid = NastiRouter_1_io_master_b_valid;
  assign io_masters_1_w_ready = NastiRouter_1_io_master_w_ready;
  assign io_masters_1_aw_ready = NastiRouter_1_io_master_aw_ready;
  NastiRouter_0 NastiRouter(.clk(clk), .reset(reset),
       .io_master_aw_ready( NastiRouter_io_master_aw_ready ),
       .io_master_aw_valid( io_masters_0_aw_valid ),
       .io_master_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_master_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_master_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_master_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_master_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_master_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_master_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_master_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_master_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_master_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_master_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_master_w_ready( NastiRouter_io_master_w_ready ),
       .io_master_w_valid( io_masters_0_w_valid ),
       .io_master_w_bits_data( io_masters_0_w_bits_data ),
       .io_master_w_bits_last( io_masters_0_w_bits_last ),
       .io_master_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_master_w_bits_user( io_masters_0_w_bits_user ),
       .io_master_b_ready( io_masters_0_b_ready ),
       .io_master_b_valid( NastiRouter_io_master_b_valid ),
       .io_master_b_bits_resp( NastiRouter_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiRouter_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiRouter_io_master_b_bits_user ),
       .io_master_ar_ready( NastiRouter_io_master_ar_ready ),
       .io_master_ar_valid( io_masters_0_ar_valid ),
       .io_master_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_master_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_master_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_master_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_master_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_master_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_master_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_master_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_master_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_master_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_master_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_master_r_ready( io_masters_0_r_ready ),
       .io_master_r_valid( NastiRouter_io_master_r_valid ),
       .io_master_r_bits_resp( NastiRouter_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiRouter_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiRouter_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiRouter_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiRouter_io_master_r_bits_user ),
       .io_slave_2_aw_ready( NastiArbiter_2_io_master_0_aw_ready ),
       .io_slave_2_aw_valid( NastiRouter_io_slave_2_aw_valid ),
       .io_slave_2_aw_bits_addr( NastiRouter_io_slave_2_aw_bits_addr ),
       .io_slave_2_aw_bits_len( NastiRouter_io_slave_2_aw_bits_len ),
       .io_slave_2_aw_bits_size( NastiRouter_io_slave_2_aw_bits_size ),
       .io_slave_2_aw_bits_burst( NastiRouter_io_slave_2_aw_bits_burst ),
       .io_slave_2_aw_bits_lock( NastiRouter_io_slave_2_aw_bits_lock ),
       .io_slave_2_aw_bits_cache( NastiRouter_io_slave_2_aw_bits_cache ),
       .io_slave_2_aw_bits_prot( NastiRouter_io_slave_2_aw_bits_prot ),
       .io_slave_2_aw_bits_qos( NastiRouter_io_slave_2_aw_bits_qos ),
       .io_slave_2_aw_bits_region( NastiRouter_io_slave_2_aw_bits_region ),
       .io_slave_2_aw_bits_id( NastiRouter_io_slave_2_aw_bits_id ),
       .io_slave_2_aw_bits_user( NastiRouter_io_slave_2_aw_bits_user ),
       .io_slave_2_w_ready( NastiArbiter_2_io_master_0_w_ready ),
       .io_slave_2_w_valid( NastiRouter_io_slave_2_w_valid ),
       .io_slave_2_w_bits_data( NastiRouter_io_slave_2_w_bits_data ),
       .io_slave_2_w_bits_last( NastiRouter_io_slave_2_w_bits_last ),
       .io_slave_2_w_bits_strb( NastiRouter_io_slave_2_w_bits_strb ),
       .io_slave_2_w_bits_user( NastiRouter_io_slave_2_w_bits_user ),
       .io_slave_2_b_ready( NastiRouter_io_slave_2_b_ready ),
       .io_slave_2_b_valid( NastiArbiter_2_io_master_0_b_valid ),
       .io_slave_2_b_bits_resp( NastiArbiter_2_io_master_0_b_bits_resp ),
       .io_slave_2_b_bits_id( NastiArbiter_2_io_master_0_b_bits_id ),
       .io_slave_2_b_bits_user( NastiArbiter_2_io_master_0_b_bits_user ),
       .io_slave_2_ar_ready( NastiArbiter_2_io_master_0_ar_ready ),
       .io_slave_2_ar_valid( NastiRouter_io_slave_2_ar_valid ),
       .io_slave_2_ar_bits_addr( NastiRouter_io_slave_2_ar_bits_addr ),
       .io_slave_2_ar_bits_len( NastiRouter_io_slave_2_ar_bits_len ),
       .io_slave_2_ar_bits_size( NastiRouter_io_slave_2_ar_bits_size ),
       .io_slave_2_ar_bits_burst( NastiRouter_io_slave_2_ar_bits_burst ),
       .io_slave_2_ar_bits_lock( NastiRouter_io_slave_2_ar_bits_lock ),
       .io_slave_2_ar_bits_cache( NastiRouter_io_slave_2_ar_bits_cache ),
       .io_slave_2_ar_bits_prot( NastiRouter_io_slave_2_ar_bits_prot ),
       .io_slave_2_ar_bits_qos( NastiRouter_io_slave_2_ar_bits_qos ),
       .io_slave_2_ar_bits_region( NastiRouter_io_slave_2_ar_bits_region ),
       .io_slave_2_ar_bits_id( NastiRouter_io_slave_2_ar_bits_id ),
       .io_slave_2_ar_bits_user( NastiRouter_io_slave_2_ar_bits_user ),
       .io_slave_2_r_ready( NastiRouter_io_slave_2_r_ready ),
       .io_slave_2_r_valid( NastiArbiter_2_io_master_0_r_valid ),
       .io_slave_2_r_bits_resp( NastiArbiter_2_io_master_0_r_bits_resp ),
       .io_slave_2_r_bits_data( NastiArbiter_2_io_master_0_r_bits_data ),
       .io_slave_2_r_bits_last( NastiArbiter_2_io_master_0_r_bits_last ),
       .io_slave_2_r_bits_id( NastiArbiter_2_io_master_0_r_bits_id ),
       .io_slave_2_r_bits_user( NastiArbiter_2_io_master_0_r_bits_user ),
       .io_slave_1_aw_ready( NastiArbiter_1_io_master_0_aw_ready ),
       .io_slave_1_aw_valid( NastiRouter_io_slave_1_aw_valid ),
       .io_slave_1_aw_bits_addr( NastiRouter_io_slave_1_aw_bits_addr ),
       .io_slave_1_aw_bits_len( NastiRouter_io_slave_1_aw_bits_len ),
       .io_slave_1_aw_bits_size( NastiRouter_io_slave_1_aw_bits_size ),
       .io_slave_1_aw_bits_burst( NastiRouter_io_slave_1_aw_bits_burst ),
       .io_slave_1_aw_bits_lock( NastiRouter_io_slave_1_aw_bits_lock ),
       .io_slave_1_aw_bits_cache( NastiRouter_io_slave_1_aw_bits_cache ),
       .io_slave_1_aw_bits_prot( NastiRouter_io_slave_1_aw_bits_prot ),
       .io_slave_1_aw_bits_qos( NastiRouter_io_slave_1_aw_bits_qos ),
       .io_slave_1_aw_bits_region( NastiRouter_io_slave_1_aw_bits_region ),
       .io_slave_1_aw_bits_id( NastiRouter_io_slave_1_aw_bits_id ),
       .io_slave_1_aw_bits_user( NastiRouter_io_slave_1_aw_bits_user ),
       .io_slave_1_w_ready( NastiArbiter_1_io_master_0_w_ready ),
       .io_slave_1_w_valid( NastiRouter_io_slave_1_w_valid ),
       .io_slave_1_w_bits_data( NastiRouter_io_slave_1_w_bits_data ),
       .io_slave_1_w_bits_last( NastiRouter_io_slave_1_w_bits_last ),
       .io_slave_1_w_bits_strb( NastiRouter_io_slave_1_w_bits_strb ),
       .io_slave_1_w_bits_user( NastiRouter_io_slave_1_w_bits_user ),
       .io_slave_1_b_ready( NastiRouter_io_slave_1_b_ready ),
       .io_slave_1_b_valid( NastiArbiter_1_io_master_0_b_valid ),
       .io_slave_1_b_bits_resp( NastiArbiter_1_io_master_0_b_bits_resp ),
       .io_slave_1_b_bits_id( NastiArbiter_1_io_master_0_b_bits_id ),
       .io_slave_1_b_bits_user( NastiArbiter_1_io_master_0_b_bits_user ),
       .io_slave_1_ar_ready( NastiArbiter_1_io_master_0_ar_ready ),
       .io_slave_1_ar_valid( NastiRouter_io_slave_1_ar_valid ),
       .io_slave_1_ar_bits_addr( NastiRouter_io_slave_1_ar_bits_addr ),
       .io_slave_1_ar_bits_len( NastiRouter_io_slave_1_ar_bits_len ),
       .io_slave_1_ar_bits_size( NastiRouter_io_slave_1_ar_bits_size ),
       .io_slave_1_ar_bits_burst( NastiRouter_io_slave_1_ar_bits_burst ),
       .io_slave_1_ar_bits_lock( NastiRouter_io_slave_1_ar_bits_lock ),
       .io_slave_1_ar_bits_cache( NastiRouter_io_slave_1_ar_bits_cache ),
       .io_slave_1_ar_bits_prot( NastiRouter_io_slave_1_ar_bits_prot ),
       .io_slave_1_ar_bits_qos( NastiRouter_io_slave_1_ar_bits_qos ),
       .io_slave_1_ar_bits_region( NastiRouter_io_slave_1_ar_bits_region ),
       .io_slave_1_ar_bits_id( NastiRouter_io_slave_1_ar_bits_id ),
       .io_slave_1_ar_bits_user( NastiRouter_io_slave_1_ar_bits_user ),
       .io_slave_1_r_ready( NastiRouter_io_slave_1_r_ready ),
       .io_slave_1_r_valid( NastiArbiter_1_io_master_0_r_valid ),
       .io_slave_1_r_bits_resp( NastiArbiter_1_io_master_0_r_bits_resp ),
       .io_slave_1_r_bits_data( NastiArbiter_1_io_master_0_r_bits_data ),
       .io_slave_1_r_bits_last( NastiArbiter_1_io_master_0_r_bits_last ),
       .io_slave_1_r_bits_id( NastiArbiter_1_io_master_0_r_bits_id ),
       .io_slave_1_r_bits_user( NastiArbiter_1_io_master_0_r_bits_user ),
       .io_slave_0_aw_ready( NastiArbiter_io_master_0_aw_ready ),
       .io_slave_0_aw_valid( NastiRouter_io_slave_0_aw_valid ),
       .io_slave_0_aw_bits_addr( NastiRouter_io_slave_0_aw_bits_addr ),
       .io_slave_0_aw_bits_len( NastiRouter_io_slave_0_aw_bits_len ),
       .io_slave_0_aw_bits_size( NastiRouter_io_slave_0_aw_bits_size ),
       .io_slave_0_aw_bits_burst( NastiRouter_io_slave_0_aw_bits_burst ),
       .io_slave_0_aw_bits_lock( NastiRouter_io_slave_0_aw_bits_lock ),
       .io_slave_0_aw_bits_cache( NastiRouter_io_slave_0_aw_bits_cache ),
       .io_slave_0_aw_bits_prot( NastiRouter_io_slave_0_aw_bits_prot ),
       .io_slave_0_aw_bits_qos( NastiRouter_io_slave_0_aw_bits_qos ),
       .io_slave_0_aw_bits_region( NastiRouter_io_slave_0_aw_bits_region ),
       .io_slave_0_aw_bits_id( NastiRouter_io_slave_0_aw_bits_id ),
       .io_slave_0_aw_bits_user( NastiRouter_io_slave_0_aw_bits_user ),
       .io_slave_0_w_ready( NastiArbiter_io_master_0_w_ready ),
       .io_slave_0_w_valid( NastiRouter_io_slave_0_w_valid ),
       .io_slave_0_w_bits_data( NastiRouter_io_slave_0_w_bits_data ),
       .io_slave_0_w_bits_last( NastiRouter_io_slave_0_w_bits_last ),
       .io_slave_0_w_bits_strb( NastiRouter_io_slave_0_w_bits_strb ),
       .io_slave_0_w_bits_user( NastiRouter_io_slave_0_w_bits_user ),
       .io_slave_0_b_ready( NastiRouter_io_slave_0_b_ready ),
       .io_slave_0_b_valid( NastiArbiter_io_master_0_b_valid ),
       .io_slave_0_b_bits_resp( NastiArbiter_io_master_0_b_bits_resp ),
       .io_slave_0_b_bits_id( NastiArbiter_io_master_0_b_bits_id ),
       .io_slave_0_b_bits_user( NastiArbiter_io_master_0_b_bits_user ),
       .io_slave_0_ar_ready( NastiArbiter_io_master_0_ar_ready ),
       .io_slave_0_ar_valid( NastiRouter_io_slave_0_ar_valid ),
       .io_slave_0_ar_bits_addr( NastiRouter_io_slave_0_ar_bits_addr ),
       .io_slave_0_ar_bits_len( NastiRouter_io_slave_0_ar_bits_len ),
       .io_slave_0_ar_bits_size( NastiRouter_io_slave_0_ar_bits_size ),
       .io_slave_0_ar_bits_burst( NastiRouter_io_slave_0_ar_bits_burst ),
       .io_slave_0_ar_bits_lock( NastiRouter_io_slave_0_ar_bits_lock ),
       .io_slave_0_ar_bits_cache( NastiRouter_io_slave_0_ar_bits_cache ),
       .io_slave_0_ar_bits_prot( NastiRouter_io_slave_0_ar_bits_prot ),
       .io_slave_0_ar_bits_qos( NastiRouter_io_slave_0_ar_bits_qos ),
       .io_slave_0_ar_bits_region( NastiRouter_io_slave_0_ar_bits_region ),
       .io_slave_0_ar_bits_id( NastiRouter_io_slave_0_ar_bits_id ),
       .io_slave_0_ar_bits_user( NastiRouter_io_slave_0_ar_bits_user ),
       .io_slave_0_r_ready( NastiRouter_io_slave_0_r_ready ),
       .io_slave_0_r_valid( NastiArbiter_io_master_0_r_valid ),
       .io_slave_0_r_bits_resp( NastiArbiter_io_master_0_r_bits_resp ),
       .io_slave_0_r_bits_data( NastiArbiter_io_master_0_r_bits_data ),
       .io_slave_0_r_bits_last( NastiArbiter_io_master_0_r_bits_last ),
       .io_slave_0_r_bits_id( NastiArbiter_io_master_0_r_bits_id ),
       .io_slave_0_r_bits_user( NastiArbiter_io_master_0_r_bits_user )
  );
  NastiRouter_0 NastiRouter_1(.clk(clk), .reset(reset),
       .io_master_aw_ready( NastiRouter_1_io_master_aw_ready ),
       .io_master_aw_valid( io_masters_1_aw_valid ),
       .io_master_aw_bits_addr( io_masters_1_aw_bits_addr ),
       .io_master_aw_bits_len( io_masters_1_aw_bits_len ),
       .io_master_aw_bits_size( io_masters_1_aw_bits_size ),
       .io_master_aw_bits_burst( io_masters_1_aw_bits_burst ),
       .io_master_aw_bits_lock( io_masters_1_aw_bits_lock ),
       .io_master_aw_bits_cache( io_masters_1_aw_bits_cache ),
       .io_master_aw_bits_prot( io_masters_1_aw_bits_prot ),
       .io_master_aw_bits_qos( io_masters_1_aw_bits_qos ),
       .io_master_aw_bits_region( io_masters_1_aw_bits_region ),
       .io_master_aw_bits_id( io_masters_1_aw_bits_id ),
       .io_master_aw_bits_user( io_masters_1_aw_bits_user ),
       .io_master_w_ready( NastiRouter_1_io_master_w_ready ),
       .io_master_w_valid( io_masters_1_w_valid ),
       .io_master_w_bits_data( io_masters_1_w_bits_data ),
       .io_master_w_bits_last( io_masters_1_w_bits_last ),
       .io_master_w_bits_strb( io_masters_1_w_bits_strb ),
       .io_master_w_bits_user( io_masters_1_w_bits_user ),
       .io_master_b_ready( io_masters_1_b_ready ),
       .io_master_b_valid( NastiRouter_1_io_master_b_valid ),
       .io_master_b_bits_resp( NastiRouter_1_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiRouter_1_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiRouter_1_io_master_b_bits_user ),
       .io_master_ar_ready( NastiRouter_1_io_master_ar_ready ),
       .io_master_ar_valid( io_masters_1_ar_valid ),
       .io_master_ar_bits_addr( io_masters_1_ar_bits_addr ),
       .io_master_ar_bits_len( io_masters_1_ar_bits_len ),
       .io_master_ar_bits_size( io_masters_1_ar_bits_size ),
       .io_master_ar_bits_burst( io_masters_1_ar_bits_burst ),
       .io_master_ar_bits_lock( io_masters_1_ar_bits_lock ),
       .io_master_ar_bits_cache( io_masters_1_ar_bits_cache ),
       .io_master_ar_bits_prot( io_masters_1_ar_bits_prot ),
       .io_master_ar_bits_qos( io_masters_1_ar_bits_qos ),
       .io_master_ar_bits_region( io_masters_1_ar_bits_region ),
       .io_master_ar_bits_id( io_masters_1_ar_bits_id ),
       .io_master_ar_bits_user( io_masters_1_ar_bits_user ),
       .io_master_r_ready( io_masters_1_r_ready ),
       .io_master_r_valid( NastiRouter_1_io_master_r_valid ),
       .io_master_r_bits_resp( NastiRouter_1_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiRouter_1_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiRouter_1_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiRouter_1_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiRouter_1_io_master_r_bits_user ),
       .io_slave_2_aw_ready( NastiArbiter_2_io_master_1_aw_ready ),
       .io_slave_2_aw_valid( NastiRouter_1_io_slave_2_aw_valid ),
       .io_slave_2_aw_bits_addr( NastiRouter_1_io_slave_2_aw_bits_addr ),
       .io_slave_2_aw_bits_len( NastiRouter_1_io_slave_2_aw_bits_len ),
       .io_slave_2_aw_bits_size( NastiRouter_1_io_slave_2_aw_bits_size ),
       .io_slave_2_aw_bits_burst( NastiRouter_1_io_slave_2_aw_bits_burst ),
       .io_slave_2_aw_bits_lock( NastiRouter_1_io_slave_2_aw_bits_lock ),
       .io_slave_2_aw_bits_cache( NastiRouter_1_io_slave_2_aw_bits_cache ),
       .io_slave_2_aw_bits_prot( NastiRouter_1_io_slave_2_aw_bits_prot ),
       .io_slave_2_aw_bits_qos( NastiRouter_1_io_slave_2_aw_bits_qos ),
       .io_slave_2_aw_bits_region( NastiRouter_1_io_slave_2_aw_bits_region ),
       .io_slave_2_aw_bits_id( NastiRouter_1_io_slave_2_aw_bits_id ),
       .io_slave_2_aw_bits_user( NastiRouter_1_io_slave_2_aw_bits_user ),
       .io_slave_2_w_ready( NastiArbiter_2_io_master_1_w_ready ),
       .io_slave_2_w_valid( NastiRouter_1_io_slave_2_w_valid ),
       .io_slave_2_w_bits_data( NastiRouter_1_io_slave_2_w_bits_data ),
       .io_slave_2_w_bits_last( NastiRouter_1_io_slave_2_w_bits_last ),
       .io_slave_2_w_bits_strb( NastiRouter_1_io_slave_2_w_bits_strb ),
       .io_slave_2_w_bits_user( NastiRouter_1_io_slave_2_w_bits_user ),
       .io_slave_2_b_ready( NastiRouter_1_io_slave_2_b_ready ),
       .io_slave_2_b_valid( NastiArbiter_2_io_master_1_b_valid ),
       .io_slave_2_b_bits_resp( NastiArbiter_2_io_master_1_b_bits_resp ),
       .io_slave_2_b_bits_id( NastiArbiter_2_io_master_1_b_bits_id ),
       .io_slave_2_b_bits_user( NastiArbiter_2_io_master_1_b_bits_user ),
       .io_slave_2_ar_ready( NastiArbiter_2_io_master_1_ar_ready ),
       .io_slave_2_ar_valid( NastiRouter_1_io_slave_2_ar_valid ),
       .io_slave_2_ar_bits_addr( NastiRouter_1_io_slave_2_ar_bits_addr ),
       .io_slave_2_ar_bits_len( NastiRouter_1_io_slave_2_ar_bits_len ),
       .io_slave_2_ar_bits_size( NastiRouter_1_io_slave_2_ar_bits_size ),
       .io_slave_2_ar_bits_burst( NastiRouter_1_io_slave_2_ar_bits_burst ),
       .io_slave_2_ar_bits_lock( NastiRouter_1_io_slave_2_ar_bits_lock ),
       .io_slave_2_ar_bits_cache( NastiRouter_1_io_slave_2_ar_bits_cache ),
       .io_slave_2_ar_bits_prot( NastiRouter_1_io_slave_2_ar_bits_prot ),
       .io_slave_2_ar_bits_qos( NastiRouter_1_io_slave_2_ar_bits_qos ),
       .io_slave_2_ar_bits_region( NastiRouter_1_io_slave_2_ar_bits_region ),
       .io_slave_2_ar_bits_id( NastiRouter_1_io_slave_2_ar_bits_id ),
       .io_slave_2_ar_bits_user( NastiRouter_1_io_slave_2_ar_bits_user ),
       .io_slave_2_r_ready( NastiRouter_1_io_slave_2_r_ready ),
       .io_slave_2_r_valid( NastiArbiter_2_io_master_1_r_valid ),
       .io_slave_2_r_bits_resp( NastiArbiter_2_io_master_1_r_bits_resp ),
       .io_slave_2_r_bits_data( NastiArbiter_2_io_master_1_r_bits_data ),
       .io_slave_2_r_bits_last( NastiArbiter_2_io_master_1_r_bits_last ),
       .io_slave_2_r_bits_id( NastiArbiter_2_io_master_1_r_bits_id ),
       .io_slave_2_r_bits_user( NastiArbiter_2_io_master_1_r_bits_user ),
       .io_slave_1_aw_ready( NastiArbiter_1_io_master_1_aw_ready ),
       .io_slave_1_aw_valid( NastiRouter_1_io_slave_1_aw_valid ),
       .io_slave_1_aw_bits_addr( NastiRouter_1_io_slave_1_aw_bits_addr ),
       .io_slave_1_aw_bits_len( NastiRouter_1_io_slave_1_aw_bits_len ),
       .io_slave_1_aw_bits_size( NastiRouter_1_io_slave_1_aw_bits_size ),
       .io_slave_1_aw_bits_burst( NastiRouter_1_io_slave_1_aw_bits_burst ),
       .io_slave_1_aw_bits_lock( NastiRouter_1_io_slave_1_aw_bits_lock ),
       .io_slave_1_aw_bits_cache( NastiRouter_1_io_slave_1_aw_bits_cache ),
       .io_slave_1_aw_bits_prot( NastiRouter_1_io_slave_1_aw_bits_prot ),
       .io_slave_1_aw_bits_qos( NastiRouter_1_io_slave_1_aw_bits_qos ),
       .io_slave_1_aw_bits_region( NastiRouter_1_io_slave_1_aw_bits_region ),
       .io_slave_1_aw_bits_id( NastiRouter_1_io_slave_1_aw_bits_id ),
       .io_slave_1_aw_bits_user( NastiRouter_1_io_slave_1_aw_bits_user ),
       .io_slave_1_w_ready( NastiArbiter_1_io_master_1_w_ready ),
       .io_slave_1_w_valid( NastiRouter_1_io_slave_1_w_valid ),
       .io_slave_1_w_bits_data( NastiRouter_1_io_slave_1_w_bits_data ),
       .io_slave_1_w_bits_last( NastiRouter_1_io_slave_1_w_bits_last ),
       .io_slave_1_w_bits_strb( NastiRouter_1_io_slave_1_w_bits_strb ),
       .io_slave_1_w_bits_user( NastiRouter_1_io_slave_1_w_bits_user ),
       .io_slave_1_b_ready( NastiRouter_1_io_slave_1_b_ready ),
       .io_slave_1_b_valid( NastiArbiter_1_io_master_1_b_valid ),
       .io_slave_1_b_bits_resp( NastiArbiter_1_io_master_1_b_bits_resp ),
       .io_slave_1_b_bits_id( NastiArbiter_1_io_master_1_b_bits_id ),
       .io_slave_1_b_bits_user( NastiArbiter_1_io_master_1_b_bits_user ),
       .io_slave_1_ar_ready( NastiArbiter_1_io_master_1_ar_ready ),
       .io_slave_1_ar_valid( NastiRouter_1_io_slave_1_ar_valid ),
       .io_slave_1_ar_bits_addr( NastiRouter_1_io_slave_1_ar_bits_addr ),
       .io_slave_1_ar_bits_len( NastiRouter_1_io_slave_1_ar_bits_len ),
       .io_slave_1_ar_bits_size( NastiRouter_1_io_slave_1_ar_bits_size ),
       .io_slave_1_ar_bits_burst( NastiRouter_1_io_slave_1_ar_bits_burst ),
       .io_slave_1_ar_bits_lock( NastiRouter_1_io_slave_1_ar_bits_lock ),
       .io_slave_1_ar_bits_cache( NastiRouter_1_io_slave_1_ar_bits_cache ),
       .io_slave_1_ar_bits_prot( NastiRouter_1_io_slave_1_ar_bits_prot ),
       .io_slave_1_ar_bits_qos( NastiRouter_1_io_slave_1_ar_bits_qos ),
       .io_slave_1_ar_bits_region( NastiRouter_1_io_slave_1_ar_bits_region ),
       .io_slave_1_ar_bits_id( NastiRouter_1_io_slave_1_ar_bits_id ),
       .io_slave_1_ar_bits_user( NastiRouter_1_io_slave_1_ar_bits_user ),
       .io_slave_1_r_ready( NastiRouter_1_io_slave_1_r_ready ),
       .io_slave_1_r_valid( NastiArbiter_1_io_master_1_r_valid ),
       .io_slave_1_r_bits_resp( NastiArbiter_1_io_master_1_r_bits_resp ),
       .io_slave_1_r_bits_data( NastiArbiter_1_io_master_1_r_bits_data ),
       .io_slave_1_r_bits_last( NastiArbiter_1_io_master_1_r_bits_last ),
       .io_slave_1_r_bits_id( NastiArbiter_1_io_master_1_r_bits_id ),
       .io_slave_1_r_bits_user( NastiArbiter_1_io_master_1_r_bits_user ),
       .io_slave_0_aw_ready( NastiArbiter_io_master_1_aw_ready ),
       .io_slave_0_aw_valid( NastiRouter_1_io_slave_0_aw_valid ),
       .io_slave_0_aw_bits_addr( NastiRouter_1_io_slave_0_aw_bits_addr ),
       .io_slave_0_aw_bits_len( NastiRouter_1_io_slave_0_aw_bits_len ),
       .io_slave_0_aw_bits_size( NastiRouter_1_io_slave_0_aw_bits_size ),
       .io_slave_0_aw_bits_burst( NastiRouter_1_io_slave_0_aw_bits_burst ),
       .io_slave_0_aw_bits_lock( NastiRouter_1_io_slave_0_aw_bits_lock ),
       .io_slave_0_aw_bits_cache( NastiRouter_1_io_slave_0_aw_bits_cache ),
       .io_slave_0_aw_bits_prot( NastiRouter_1_io_slave_0_aw_bits_prot ),
       .io_slave_0_aw_bits_qos( NastiRouter_1_io_slave_0_aw_bits_qos ),
       .io_slave_0_aw_bits_region( NastiRouter_1_io_slave_0_aw_bits_region ),
       .io_slave_0_aw_bits_id( NastiRouter_1_io_slave_0_aw_bits_id ),
       .io_slave_0_aw_bits_user( NastiRouter_1_io_slave_0_aw_bits_user ),
       .io_slave_0_w_ready( NastiArbiter_io_master_1_w_ready ),
       .io_slave_0_w_valid( NastiRouter_1_io_slave_0_w_valid ),
       .io_slave_0_w_bits_data( NastiRouter_1_io_slave_0_w_bits_data ),
       .io_slave_0_w_bits_last( NastiRouter_1_io_slave_0_w_bits_last ),
       .io_slave_0_w_bits_strb( NastiRouter_1_io_slave_0_w_bits_strb ),
       .io_slave_0_w_bits_user( NastiRouter_1_io_slave_0_w_bits_user ),
       .io_slave_0_b_ready( NastiRouter_1_io_slave_0_b_ready ),
       .io_slave_0_b_valid( NastiArbiter_io_master_1_b_valid ),
       .io_slave_0_b_bits_resp( NastiArbiter_io_master_1_b_bits_resp ),
       .io_slave_0_b_bits_id( NastiArbiter_io_master_1_b_bits_id ),
       .io_slave_0_b_bits_user( NastiArbiter_io_master_1_b_bits_user ),
       .io_slave_0_ar_ready( NastiArbiter_io_master_1_ar_ready ),
       .io_slave_0_ar_valid( NastiRouter_1_io_slave_0_ar_valid ),
       .io_slave_0_ar_bits_addr( NastiRouter_1_io_slave_0_ar_bits_addr ),
       .io_slave_0_ar_bits_len( NastiRouter_1_io_slave_0_ar_bits_len ),
       .io_slave_0_ar_bits_size( NastiRouter_1_io_slave_0_ar_bits_size ),
       .io_slave_0_ar_bits_burst( NastiRouter_1_io_slave_0_ar_bits_burst ),
       .io_slave_0_ar_bits_lock( NastiRouter_1_io_slave_0_ar_bits_lock ),
       .io_slave_0_ar_bits_cache( NastiRouter_1_io_slave_0_ar_bits_cache ),
       .io_slave_0_ar_bits_prot( NastiRouter_1_io_slave_0_ar_bits_prot ),
       .io_slave_0_ar_bits_qos( NastiRouter_1_io_slave_0_ar_bits_qos ),
       .io_slave_0_ar_bits_region( NastiRouter_1_io_slave_0_ar_bits_region ),
       .io_slave_0_ar_bits_id( NastiRouter_1_io_slave_0_ar_bits_id ),
       .io_slave_0_ar_bits_user( NastiRouter_1_io_slave_0_ar_bits_user ),
       .io_slave_0_r_ready( NastiRouter_1_io_slave_0_r_ready ),
       .io_slave_0_r_valid( NastiArbiter_io_master_1_r_valid ),
       .io_slave_0_r_bits_resp( NastiArbiter_io_master_1_r_bits_resp ),
       .io_slave_0_r_bits_data( NastiArbiter_io_master_1_r_bits_data ),
       .io_slave_0_r_bits_last( NastiArbiter_io_master_1_r_bits_last ),
       .io_slave_0_r_bits_id( NastiArbiter_io_master_1_r_bits_id ),
       .io_slave_0_r_bits_user( NastiArbiter_io_master_1_r_bits_user )
  );
  NastiArbiter NastiArbiter(.clk(clk), .reset(reset),
       .io_master_1_aw_ready( NastiArbiter_io_master_1_aw_ready ),
       .io_master_1_aw_valid( NastiRouter_1_io_slave_0_aw_valid ),
       .io_master_1_aw_bits_addr( NastiRouter_1_io_slave_0_aw_bits_addr ),
       .io_master_1_aw_bits_len( NastiRouter_1_io_slave_0_aw_bits_len ),
       .io_master_1_aw_bits_size( NastiRouter_1_io_slave_0_aw_bits_size ),
       .io_master_1_aw_bits_burst( NastiRouter_1_io_slave_0_aw_bits_burst ),
       .io_master_1_aw_bits_lock( NastiRouter_1_io_slave_0_aw_bits_lock ),
       .io_master_1_aw_bits_cache( NastiRouter_1_io_slave_0_aw_bits_cache ),
       .io_master_1_aw_bits_prot( NastiRouter_1_io_slave_0_aw_bits_prot ),
       .io_master_1_aw_bits_qos( NastiRouter_1_io_slave_0_aw_bits_qos ),
       .io_master_1_aw_bits_region( NastiRouter_1_io_slave_0_aw_bits_region ),
       .io_master_1_aw_bits_id( NastiRouter_1_io_slave_0_aw_bits_id ),
       .io_master_1_aw_bits_user( NastiRouter_1_io_slave_0_aw_bits_user ),
       .io_master_1_w_ready( NastiArbiter_io_master_1_w_ready ),
       .io_master_1_w_valid( NastiRouter_1_io_slave_0_w_valid ),
       .io_master_1_w_bits_data( NastiRouter_1_io_slave_0_w_bits_data ),
       .io_master_1_w_bits_last( NastiRouter_1_io_slave_0_w_bits_last ),
       .io_master_1_w_bits_strb( NastiRouter_1_io_slave_0_w_bits_strb ),
       .io_master_1_w_bits_user( NastiRouter_1_io_slave_0_w_bits_user ),
       .io_master_1_b_ready( NastiRouter_1_io_slave_0_b_ready ),
       .io_master_1_b_valid( NastiArbiter_io_master_1_b_valid ),
       .io_master_1_b_bits_resp( NastiArbiter_io_master_1_b_bits_resp ),
       .io_master_1_b_bits_id( NastiArbiter_io_master_1_b_bits_id ),
       .io_master_1_b_bits_user( NastiArbiter_io_master_1_b_bits_user ),
       .io_master_1_ar_ready( NastiArbiter_io_master_1_ar_ready ),
       .io_master_1_ar_valid( NastiRouter_1_io_slave_0_ar_valid ),
       .io_master_1_ar_bits_addr( NastiRouter_1_io_slave_0_ar_bits_addr ),
       .io_master_1_ar_bits_len( NastiRouter_1_io_slave_0_ar_bits_len ),
       .io_master_1_ar_bits_size( NastiRouter_1_io_slave_0_ar_bits_size ),
       .io_master_1_ar_bits_burst( NastiRouter_1_io_slave_0_ar_bits_burst ),
       .io_master_1_ar_bits_lock( NastiRouter_1_io_slave_0_ar_bits_lock ),
       .io_master_1_ar_bits_cache( NastiRouter_1_io_slave_0_ar_bits_cache ),
       .io_master_1_ar_bits_prot( NastiRouter_1_io_slave_0_ar_bits_prot ),
       .io_master_1_ar_bits_qos( NastiRouter_1_io_slave_0_ar_bits_qos ),
       .io_master_1_ar_bits_region( NastiRouter_1_io_slave_0_ar_bits_region ),
       .io_master_1_ar_bits_id( NastiRouter_1_io_slave_0_ar_bits_id ),
       .io_master_1_ar_bits_user( NastiRouter_1_io_slave_0_ar_bits_user ),
       .io_master_1_r_ready( NastiRouter_1_io_slave_0_r_ready ),
       .io_master_1_r_valid( NastiArbiter_io_master_1_r_valid ),
       .io_master_1_r_bits_resp( NastiArbiter_io_master_1_r_bits_resp ),
       .io_master_1_r_bits_data( NastiArbiter_io_master_1_r_bits_data ),
       .io_master_1_r_bits_last( NastiArbiter_io_master_1_r_bits_last ),
       .io_master_1_r_bits_id( NastiArbiter_io_master_1_r_bits_id ),
       .io_master_1_r_bits_user( NastiArbiter_io_master_1_r_bits_user ),
       .io_master_0_aw_ready( NastiArbiter_io_master_0_aw_ready ),
       .io_master_0_aw_valid( NastiRouter_io_slave_0_aw_valid ),
       .io_master_0_aw_bits_addr( NastiRouter_io_slave_0_aw_bits_addr ),
       .io_master_0_aw_bits_len( NastiRouter_io_slave_0_aw_bits_len ),
       .io_master_0_aw_bits_size( NastiRouter_io_slave_0_aw_bits_size ),
       .io_master_0_aw_bits_burst( NastiRouter_io_slave_0_aw_bits_burst ),
       .io_master_0_aw_bits_lock( NastiRouter_io_slave_0_aw_bits_lock ),
       .io_master_0_aw_bits_cache( NastiRouter_io_slave_0_aw_bits_cache ),
       .io_master_0_aw_bits_prot( NastiRouter_io_slave_0_aw_bits_prot ),
       .io_master_0_aw_bits_qos( NastiRouter_io_slave_0_aw_bits_qos ),
       .io_master_0_aw_bits_region( NastiRouter_io_slave_0_aw_bits_region ),
       .io_master_0_aw_bits_id( NastiRouter_io_slave_0_aw_bits_id ),
       .io_master_0_aw_bits_user( NastiRouter_io_slave_0_aw_bits_user ),
       .io_master_0_w_ready( NastiArbiter_io_master_0_w_ready ),
       .io_master_0_w_valid( NastiRouter_io_slave_0_w_valid ),
       .io_master_0_w_bits_data( NastiRouter_io_slave_0_w_bits_data ),
       .io_master_0_w_bits_last( NastiRouter_io_slave_0_w_bits_last ),
       .io_master_0_w_bits_strb( NastiRouter_io_slave_0_w_bits_strb ),
       .io_master_0_w_bits_user( NastiRouter_io_slave_0_w_bits_user ),
       .io_master_0_b_ready( NastiRouter_io_slave_0_b_ready ),
       .io_master_0_b_valid( NastiArbiter_io_master_0_b_valid ),
       .io_master_0_b_bits_resp( NastiArbiter_io_master_0_b_bits_resp ),
       .io_master_0_b_bits_id( NastiArbiter_io_master_0_b_bits_id ),
       .io_master_0_b_bits_user( NastiArbiter_io_master_0_b_bits_user ),
       .io_master_0_ar_ready( NastiArbiter_io_master_0_ar_ready ),
       .io_master_0_ar_valid( NastiRouter_io_slave_0_ar_valid ),
       .io_master_0_ar_bits_addr( NastiRouter_io_slave_0_ar_bits_addr ),
       .io_master_0_ar_bits_len( NastiRouter_io_slave_0_ar_bits_len ),
       .io_master_0_ar_bits_size( NastiRouter_io_slave_0_ar_bits_size ),
       .io_master_0_ar_bits_burst( NastiRouter_io_slave_0_ar_bits_burst ),
       .io_master_0_ar_bits_lock( NastiRouter_io_slave_0_ar_bits_lock ),
       .io_master_0_ar_bits_cache( NastiRouter_io_slave_0_ar_bits_cache ),
       .io_master_0_ar_bits_prot( NastiRouter_io_slave_0_ar_bits_prot ),
       .io_master_0_ar_bits_qos( NastiRouter_io_slave_0_ar_bits_qos ),
       .io_master_0_ar_bits_region( NastiRouter_io_slave_0_ar_bits_region ),
       .io_master_0_ar_bits_id( NastiRouter_io_slave_0_ar_bits_id ),
       .io_master_0_ar_bits_user( NastiRouter_io_slave_0_ar_bits_user ),
       .io_master_0_r_ready( NastiRouter_io_slave_0_r_ready ),
       .io_master_0_r_valid( NastiArbiter_io_master_0_r_valid ),
       .io_master_0_r_bits_resp( NastiArbiter_io_master_0_r_bits_resp ),
       .io_master_0_r_bits_data( NastiArbiter_io_master_0_r_bits_data ),
       .io_master_0_r_bits_last( NastiArbiter_io_master_0_r_bits_last ),
       .io_master_0_r_bits_id( NastiArbiter_io_master_0_r_bits_id ),
       .io_master_0_r_bits_user( NastiArbiter_io_master_0_r_bits_user ),
       .io_slave_aw_ready( io_slaves_0_aw_ready ),
       .io_slave_aw_valid( NastiArbiter_io_slave_aw_valid ),
       .io_slave_aw_bits_addr( NastiArbiter_io_slave_aw_bits_addr ),
       .io_slave_aw_bits_len( NastiArbiter_io_slave_aw_bits_len ),
       .io_slave_aw_bits_size( NastiArbiter_io_slave_aw_bits_size ),
       .io_slave_aw_bits_burst( NastiArbiter_io_slave_aw_bits_burst ),
       .io_slave_aw_bits_lock( NastiArbiter_io_slave_aw_bits_lock ),
       .io_slave_aw_bits_cache( NastiArbiter_io_slave_aw_bits_cache ),
       .io_slave_aw_bits_prot( NastiArbiter_io_slave_aw_bits_prot ),
       .io_slave_aw_bits_qos( NastiArbiter_io_slave_aw_bits_qos ),
       .io_slave_aw_bits_region( NastiArbiter_io_slave_aw_bits_region ),
       .io_slave_aw_bits_id( NastiArbiter_io_slave_aw_bits_id ),
       .io_slave_aw_bits_user( NastiArbiter_io_slave_aw_bits_user ),
       .io_slave_w_ready( io_slaves_0_w_ready ),
       .io_slave_w_valid( NastiArbiter_io_slave_w_valid ),
       .io_slave_w_bits_data( NastiArbiter_io_slave_w_bits_data ),
       .io_slave_w_bits_last( NastiArbiter_io_slave_w_bits_last ),
       .io_slave_w_bits_strb( NastiArbiter_io_slave_w_bits_strb ),
       .io_slave_w_bits_user( NastiArbiter_io_slave_w_bits_user ),
       .io_slave_b_ready( NastiArbiter_io_slave_b_ready ),
       .io_slave_b_valid( io_slaves_0_b_valid ),
       .io_slave_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slave_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slave_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slave_ar_ready( io_slaves_0_ar_ready ),
       .io_slave_ar_valid( NastiArbiter_io_slave_ar_valid ),
       .io_slave_ar_bits_addr( NastiArbiter_io_slave_ar_bits_addr ),
       .io_slave_ar_bits_len( NastiArbiter_io_slave_ar_bits_len ),
       .io_slave_ar_bits_size( NastiArbiter_io_slave_ar_bits_size ),
       .io_slave_ar_bits_burst( NastiArbiter_io_slave_ar_bits_burst ),
       .io_slave_ar_bits_lock( NastiArbiter_io_slave_ar_bits_lock ),
       .io_slave_ar_bits_cache( NastiArbiter_io_slave_ar_bits_cache ),
       .io_slave_ar_bits_prot( NastiArbiter_io_slave_ar_bits_prot ),
       .io_slave_ar_bits_qos( NastiArbiter_io_slave_ar_bits_qos ),
       .io_slave_ar_bits_region( NastiArbiter_io_slave_ar_bits_region ),
       .io_slave_ar_bits_id( NastiArbiter_io_slave_ar_bits_id ),
       .io_slave_ar_bits_user( NastiArbiter_io_slave_ar_bits_user ),
       .io_slave_r_ready( NastiArbiter_io_slave_r_ready ),
       .io_slave_r_valid( io_slaves_0_r_valid ),
       .io_slave_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slave_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slave_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slave_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slave_r_bits_user( io_slaves_0_r_bits_user )
  );
  NastiArbiter NastiArbiter_1(.clk(clk), .reset(reset),
       .io_master_1_aw_ready( NastiArbiter_1_io_master_1_aw_ready ),
       .io_master_1_aw_valid( NastiRouter_1_io_slave_1_aw_valid ),
       .io_master_1_aw_bits_addr( NastiRouter_1_io_slave_1_aw_bits_addr ),
       .io_master_1_aw_bits_len( NastiRouter_1_io_slave_1_aw_bits_len ),
       .io_master_1_aw_bits_size( NastiRouter_1_io_slave_1_aw_bits_size ),
       .io_master_1_aw_bits_burst( NastiRouter_1_io_slave_1_aw_bits_burst ),
       .io_master_1_aw_bits_lock( NastiRouter_1_io_slave_1_aw_bits_lock ),
       .io_master_1_aw_bits_cache( NastiRouter_1_io_slave_1_aw_bits_cache ),
       .io_master_1_aw_bits_prot( NastiRouter_1_io_slave_1_aw_bits_prot ),
       .io_master_1_aw_bits_qos( NastiRouter_1_io_slave_1_aw_bits_qos ),
       .io_master_1_aw_bits_region( NastiRouter_1_io_slave_1_aw_bits_region ),
       .io_master_1_aw_bits_id( NastiRouter_1_io_slave_1_aw_bits_id ),
       .io_master_1_aw_bits_user( NastiRouter_1_io_slave_1_aw_bits_user ),
       .io_master_1_w_ready( NastiArbiter_1_io_master_1_w_ready ),
       .io_master_1_w_valid( NastiRouter_1_io_slave_1_w_valid ),
       .io_master_1_w_bits_data( NastiRouter_1_io_slave_1_w_bits_data ),
       .io_master_1_w_bits_last( NastiRouter_1_io_slave_1_w_bits_last ),
       .io_master_1_w_bits_strb( NastiRouter_1_io_slave_1_w_bits_strb ),
       .io_master_1_w_bits_user( NastiRouter_1_io_slave_1_w_bits_user ),
       .io_master_1_b_ready( NastiRouter_1_io_slave_1_b_ready ),
       .io_master_1_b_valid( NastiArbiter_1_io_master_1_b_valid ),
       .io_master_1_b_bits_resp( NastiArbiter_1_io_master_1_b_bits_resp ),
       .io_master_1_b_bits_id( NastiArbiter_1_io_master_1_b_bits_id ),
       .io_master_1_b_bits_user( NastiArbiter_1_io_master_1_b_bits_user ),
       .io_master_1_ar_ready( NastiArbiter_1_io_master_1_ar_ready ),
       .io_master_1_ar_valid( NastiRouter_1_io_slave_1_ar_valid ),
       .io_master_1_ar_bits_addr( NastiRouter_1_io_slave_1_ar_bits_addr ),
       .io_master_1_ar_bits_len( NastiRouter_1_io_slave_1_ar_bits_len ),
       .io_master_1_ar_bits_size( NastiRouter_1_io_slave_1_ar_bits_size ),
       .io_master_1_ar_bits_burst( NastiRouter_1_io_slave_1_ar_bits_burst ),
       .io_master_1_ar_bits_lock( NastiRouter_1_io_slave_1_ar_bits_lock ),
       .io_master_1_ar_bits_cache( NastiRouter_1_io_slave_1_ar_bits_cache ),
       .io_master_1_ar_bits_prot( NastiRouter_1_io_slave_1_ar_bits_prot ),
       .io_master_1_ar_bits_qos( NastiRouter_1_io_slave_1_ar_bits_qos ),
       .io_master_1_ar_bits_region( NastiRouter_1_io_slave_1_ar_bits_region ),
       .io_master_1_ar_bits_id( NastiRouter_1_io_slave_1_ar_bits_id ),
       .io_master_1_ar_bits_user( NastiRouter_1_io_slave_1_ar_bits_user ),
       .io_master_1_r_ready( NastiRouter_1_io_slave_1_r_ready ),
       .io_master_1_r_valid( NastiArbiter_1_io_master_1_r_valid ),
       .io_master_1_r_bits_resp( NastiArbiter_1_io_master_1_r_bits_resp ),
       .io_master_1_r_bits_data( NastiArbiter_1_io_master_1_r_bits_data ),
       .io_master_1_r_bits_last( NastiArbiter_1_io_master_1_r_bits_last ),
       .io_master_1_r_bits_id( NastiArbiter_1_io_master_1_r_bits_id ),
       .io_master_1_r_bits_user( NastiArbiter_1_io_master_1_r_bits_user ),
       .io_master_0_aw_ready( NastiArbiter_1_io_master_0_aw_ready ),
       .io_master_0_aw_valid( NastiRouter_io_slave_1_aw_valid ),
       .io_master_0_aw_bits_addr( NastiRouter_io_slave_1_aw_bits_addr ),
       .io_master_0_aw_bits_len( NastiRouter_io_slave_1_aw_bits_len ),
       .io_master_0_aw_bits_size( NastiRouter_io_slave_1_aw_bits_size ),
       .io_master_0_aw_bits_burst( NastiRouter_io_slave_1_aw_bits_burst ),
       .io_master_0_aw_bits_lock( NastiRouter_io_slave_1_aw_bits_lock ),
       .io_master_0_aw_bits_cache( NastiRouter_io_slave_1_aw_bits_cache ),
       .io_master_0_aw_bits_prot( NastiRouter_io_slave_1_aw_bits_prot ),
       .io_master_0_aw_bits_qos( NastiRouter_io_slave_1_aw_bits_qos ),
       .io_master_0_aw_bits_region( NastiRouter_io_slave_1_aw_bits_region ),
       .io_master_0_aw_bits_id( NastiRouter_io_slave_1_aw_bits_id ),
       .io_master_0_aw_bits_user( NastiRouter_io_slave_1_aw_bits_user ),
       .io_master_0_w_ready( NastiArbiter_1_io_master_0_w_ready ),
       .io_master_0_w_valid( NastiRouter_io_slave_1_w_valid ),
       .io_master_0_w_bits_data( NastiRouter_io_slave_1_w_bits_data ),
       .io_master_0_w_bits_last( NastiRouter_io_slave_1_w_bits_last ),
       .io_master_0_w_bits_strb( NastiRouter_io_slave_1_w_bits_strb ),
       .io_master_0_w_bits_user( NastiRouter_io_slave_1_w_bits_user ),
       .io_master_0_b_ready( NastiRouter_io_slave_1_b_ready ),
       .io_master_0_b_valid( NastiArbiter_1_io_master_0_b_valid ),
       .io_master_0_b_bits_resp( NastiArbiter_1_io_master_0_b_bits_resp ),
       .io_master_0_b_bits_id( NastiArbiter_1_io_master_0_b_bits_id ),
       .io_master_0_b_bits_user( NastiArbiter_1_io_master_0_b_bits_user ),
       .io_master_0_ar_ready( NastiArbiter_1_io_master_0_ar_ready ),
       .io_master_0_ar_valid( NastiRouter_io_slave_1_ar_valid ),
       .io_master_0_ar_bits_addr( NastiRouter_io_slave_1_ar_bits_addr ),
       .io_master_0_ar_bits_len( NastiRouter_io_slave_1_ar_bits_len ),
       .io_master_0_ar_bits_size( NastiRouter_io_slave_1_ar_bits_size ),
       .io_master_0_ar_bits_burst( NastiRouter_io_slave_1_ar_bits_burst ),
       .io_master_0_ar_bits_lock( NastiRouter_io_slave_1_ar_bits_lock ),
       .io_master_0_ar_bits_cache( NastiRouter_io_slave_1_ar_bits_cache ),
       .io_master_0_ar_bits_prot( NastiRouter_io_slave_1_ar_bits_prot ),
       .io_master_0_ar_bits_qos( NastiRouter_io_slave_1_ar_bits_qos ),
       .io_master_0_ar_bits_region( NastiRouter_io_slave_1_ar_bits_region ),
       .io_master_0_ar_bits_id( NastiRouter_io_slave_1_ar_bits_id ),
       .io_master_0_ar_bits_user( NastiRouter_io_slave_1_ar_bits_user ),
       .io_master_0_r_ready( NastiRouter_io_slave_1_r_ready ),
       .io_master_0_r_valid( NastiArbiter_1_io_master_0_r_valid ),
       .io_master_0_r_bits_resp( NastiArbiter_1_io_master_0_r_bits_resp ),
       .io_master_0_r_bits_data( NastiArbiter_1_io_master_0_r_bits_data ),
       .io_master_0_r_bits_last( NastiArbiter_1_io_master_0_r_bits_last ),
       .io_master_0_r_bits_id( NastiArbiter_1_io_master_0_r_bits_id ),
       .io_master_0_r_bits_user( NastiArbiter_1_io_master_0_r_bits_user ),
       .io_slave_aw_ready( io_slaves_1_aw_ready ),
       .io_slave_aw_valid( NastiArbiter_1_io_slave_aw_valid ),
       .io_slave_aw_bits_addr( NastiArbiter_1_io_slave_aw_bits_addr ),
       .io_slave_aw_bits_len( NastiArbiter_1_io_slave_aw_bits_len ),
       .io_slave_aw_bits_size( NastiArbiter_1_io_slave_aw_bits_size ),
       .io_slave_aw_bits_burst( NastiArbiter_1_io_slave_aw_bits_burst ),
       .io_slave_aw_bits_lock( NastiArbiter_1_io_slave_aw_bits_lock ),
       .io_slave_aw_bits_cache( NastiArbiter_1_io_slave_aw_bits_cache ),
       .io_slave_aw_bits_prot( NastiArbiter_1_io_slave_aw_bits_prot ),
       .io_slave_aw_bits_qos( NastiArbiter_1_io_slave_aw_bits_qos ),
       .io_slave_aw_bits_region( NastiArbiter_1_io_slave_aw_bits_region ),
       .io_slave_aw_bits_id( NastiArbiter_1_io_slave_aw_bits_id ),
       .io_slave_aw_bits_user( NastiArbiter_1_io_slave_aw_bits_user ),
       .io_slave_w_ready( io_slaves_1_w_ready ),
       .io_slave_w_valid( NastiArbiter_1_io_slave_w_valid ),
       .io_slave_w_bits_data( NastiArbiter_1_io_slave_w_bits_data ),
       .io_slave_w_bits_last( NastiArbiter_1_io_slave_w_bits_last ),
       .io_slave_w_bits_strb( NastiArbiter_1_io_slave_w_bits_strb ),
       .io_slave_w_bits_user( NastiArbiter_1_io_slave_w_bits_user ),
       .io_slave_b_ready( NastiArbiter_1_io_slave_b_ready ),
       .io_slave_b_valid( io_slaves_1_b_valid ),
       .io_slave_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slave_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slave_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slave_ar_ready( io_slaves_1_ar_ready ),
       .io_slave_ar_valid( NastiArbiter_1_io_slave_ar_valid ),
       .io_slave_ar_bits_addr( NastiArbiter_1_io_slave_ar_bits_addr ),
       .io_slave_ar_bits_len( NastiArbiter_1_io_slave_ar_bits_len ),
       .io_slave_ar_bits_size( NastiArbiter_1_io_slave_ar_bits_size ),
       .io_slave_ar_bits_burst( NastiArbiter_1_io_slave_ar_bits_burst ),
       .io_slave_ar_bits_lock( NastiArbiter_1_io_slave_ar_bits_lock ),
       .io_slave_ar_bits_cache( NastiArbiter_1_io_slave_ar_bits_cache ),
       .io_slave_ar_bits_prot( NastiArbiter_1_io_slave_ar_bits_prot ),
       .io_slave_ar_bits_qos( NastiArbiter_1_io_slave_ar_bits_qos ),
       .io_slave_ar_bits_region( NastiArbiter_1_io_slave_ar_bits_region ),
       .io_slave_ar_bits_id( NastiArbiter_1_io_slave_ar_bits_id ),
       .io_slave_ar_bits_user( NastiArbiter_1_io_slave_ar_bits_user ),
       .io_slave_r_ready( NastiArbiter_1_io_slave_r_ready ),
       .io_slave_r_valid( io_slaves_1_r_valid ),
       .io_slave_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slave_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slave_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slave_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slave_r_bits_user( io_slaves_1_r_bits_user )
  );
  NastiArbiter NastiArbiter_2(.clk(clk), .reset(reset),
       .io_master_1_aw_ready( NastiArbiter_2_io_master_1_aw_ready ),
       .io_master_1_aw_valid( NastiRouter_1_io_slave_2_aw_valid ),
       .io_master_1_aw_bits_addr( NastiRouter_1_io_slave_2_aw_bits_addr ),
       .io_master_1_aw_bits_len( NastiRouter_1_io_slave_2_aw_bits_len ),
       .io_master_1_aw_bits_size( NastiRouter_1_io_slave_2_aw_bits_size ),
       .io_master_1_aw_bits_burst( NastiRouter_1_io_slave_2_aw_bits_burst ),
       .io_master_1_aw_bits_lock( NastiRouter_1_io_slave_2_aw_bits_lock ),
       .io_master_1_aw_bits_cache( NastiRouter_1_io_slave_2_aw_bits_cache ),
       .io_master_1_aw_bits_prot( NastiRouter_1_io_slave_2_aw_bits_prot ),
       .io_master_1_aw_bits_qos( NastiRouter_1_io_slave_2_aw_bits_qos ),
       .io_master_1_aw_bits_region( NastiRouter_1_io_slave_2_aw_bits_region ),
       .io_master_1_aw_bits_id( NastiRouter_1_io_slave_2_aw_bits_id ),
       .io_master_1_aw_bits_user( NastiRouter_1_io_slave_2_aw_bits_user ),
       .io_master_1_w_ready( NastiArbiter_2_io_master_1_w_ready ),
       .io_master_1_w_valid( NastiRouter_1_io_slave_2_w_valid ),
       .io_master_1_w_bits_data( NastiRouter_1_io_slave_2_w_bits_data ),
       .io_master_1_w_bits_last( NastiRouter_1_io_slave_2_w_bits_last ),
       .io_master_1_w_bits_strb( NastiRouter_1_io_slave_2_w_bits_strb ),
       .io_master_1_w_bits_user( NastiRouter_1_io_slave_2_w_bits_user ),
       .io_master_1_b_ready( NastiRouter_1_io_slave_2_b_ready ),
       .io_master_1_b_valid( NastiArbiter_2_io_master_1_b_valid ),
       .io_master_1_b_bits_resp( NastiArbiter_2_io_master_1_b_bits_resp ),
       .io_master_1_b_bits_id( NastiArbiter_2_io_master_1_b_bits_id ),
       .io_master_1_b_bits_user( NastiArbiter_2_io_master_1_b_bits_user ),
       .io_master_1_ar_ready( NastiArbiter_2_io_master_1_ar_ready ),
       .io_master_1_ar_valid( NastiRouter_1_io_slave_2_ar_valid ),
       .io_master_1_ar_bits_addr( NastiRouter_1_io_slave_2_ar_bits_addr ),
       .io_master_1_ar_bits_len( NastiRouter_1_io_slave_2_ar_bits_len ),
       .io_master_1_ar_bits_size( NastiRouter_1_io_slave_2_ar_bits_size ),
       .io_master_1_ar_bits_burst( NastiRouter_1_io_slave_2_ar_bits_burst ),
       .io_master_1_ar_bits_lock( NastiRouter_1_io_slave_2_ar_bits_lock ),
       .io_master_1_ar_bits_cache( NastiRouter_1_io_slave_2_ar_bits_cache ),
       .io_master_1_ar_bits_prot( NastiRouter_1_io_slave_2_ar_bits_prot ),
       .io_master_1_ar_bits_qos( NastiRouter_1_io_slave_2_ar_bits_qos ),
       .io_master_1_ar_bits_region( NastiRouter_1_io_slave_2_ar_bits_region ),
       .io_master_1_ar_bits_id( NastiRouter_1_io_slave_2_ar_bits_id ),
       .io_master_1_ar_bits_user( NastiRouter_1_io_slave_2_ar_bits_user ),
       .io_master_1_r_ready( NastiRouter_1_io_slave_2_r_ready ),
       .io_master_1_r_valid( NastiArbiter_2_io_master_1_r_valid ),
       .io_master_1_r_bits_resp( NastiArbiter_2_io_master_1_r_bits_resp ),
       .io_master_1_r_bits_data( NastiArbiter_2_io_master_1_r_bits_data ),
       .io_master_1_r_bits_last( NastiArbiter_2_io_master_1_r_bits_last ),
       .io_master_1_r_bits_id( NastiArbiter_2_io_master_1_r_bits_id ),
       .io_master_1_r_bits_user( NastiArbiter_2_io_master_1_r_bits_user ),
       .io_master_0_aw_ready( NastiArbiter_2_io_master_0_aw_ready ),
       .io_master_0_aw_valid( NastiRouter_io_slave_2_aw_valid ),
       .io_master_0_aw_bits_addr( NastiRouter_io_slave_2_aw_bits_addr ),
       .io_master_0_aw_bits_len( NastiRouter_io_slave_2_aw_bits_len ),
       .io_master_0_aw_bits_size( NastiRouter_io_slave_2_aw_bits_size ),
       .io_master_0_aw_bits_burst( NastiRouter_io_slave_2_aw_bits_burst ),
       .io_master_0_aw_bits_lock( NastiRouter_io_slave_2_aw_bits_lock ),
       .io_master_0_aw_bits_cache( NastiRouter_io_slave_2_aw_bits_cache ),
       .io_master_0_aw_bits_prot( NastiRouter_io_slave_2_aw_bits_prot ),
       .io_master_0_aw_bits_qos( NastiRouter_io_slave_2_aw_bits_qos ),
       .io_master_0_aw_bits_region( NastiRouter_io_slave_2_aw_bits_region ),
       .io_master_0_aw_bits_id( NastiRouter_io_slave_2_aw_bits_id ),
       .io_master_0_aw_bits_user( NastiRouter_io_slave_2_aw_bits_user ),
       .io_master_0_w_ready( NastiArbiter_2_io_master_0_w_ready ),
       .io_master_0_w_valid( NastiRouter_io_slave_2_w_valid ),
       .io_master_0_w_bits_data( NastiRouter_io_slave_2_w_bits_data ),
       .io_master_0_w_bits_last( NastiRouter_io_slave_2_w_bits_last ),
       .io_master_0_w_bits_strb( NastiRouter_io_slave_2_w_bits_strb ),
       .io_master_0_w_bits_user( NastiRouter_io_slave_2_w_bits_user ),
       .io_master_0_b_ready( NastiRouter_io_slave_2_b_ready ),
       .io_master_0_b_valid( NastiArbiter_2_io_master_0_b_valid ),
       .io_master_0_b_bits_resp( NastiArbiter_2_io_master_0_b_bits_resp ),
       .io_master_0_b_bits_id( NastiArbiter_2_io_master_0_b_bits_id ),
       .io_master_0_b_bits_user( NastiArbiter_2_io_master_0_b_bits_user ),
       .io_master_0_ar_ready( NastiArbiter_2_io_master_0_ar_ready ),
       .io_master_0_ar_valid( NastiRouter_io_slave_2_ar_valid ),
       .io_master_0_ar_bits_addr( NastiRouter_io_slave_2_ar_bits_addr ),
       .io_master_0_ar_bits_len( NastiRouter_io_slave_2_ar_bits_len ),
       .io_master_0_ar_bits_size( NastiRouter_io_slave_2_ar_bits_size ),
       .io_master_0_ar_bits_burst( NastiRouter_io_slave_2_ar_bits_burst ),
       .io_master_0_ar_bits_lock( NastiRouter_io_slave_2_ar_bits_lock ),
       .io_master_0_ar_bits_cache( NastiRouter_io_slave_2_ar_bits_cache ),
       .io_master_0_ar_bits_prot( NastiRouter_io_slave_2_ar_bits_prot ),
       .io_master_0_ar_bits_qos( NastiRouter_io_slave_2_ar_bits_qos ),
       .io_master_0_ar_bits_region( NastiRouter_io_slave_2_ar_bits_region ),
       .io_master_0_ar_bits_id( NastiRouter_io_slave_2_ar_bits_id ),
       .io_master_0_ar_bits_user( NastiRouter_io_slave_2_ar_bits_user ),
       .io_master_0_r_ready( NastiRouter_io_slave_2_r_ready ),
       .io_master_0_r_valid( NastiArbiter_2_io_master_0_r_valid ),
       .io_master_0_r_bits_resp( NastiArbiter_2_io_master_0_r_bits_resp ),
       .io_master_0_r_bits_data( NastiArbiter_2_io_master_0_r_bits_data ),
       .io_master_0_r_bits_last( NastiArbiter_2_io_master_0_r_bits_last ),
       .io_master_0_r_bits_id( NastiArbiter_2_io_master_0_r_bits_id ),
       .io_master_0_r_bits_user( NastiArbiter_2_io_master_0_r_bits_user ),
       .io_slave_aw_ready( io_slaves_2_aw_ready ),
       .io_slave_aw_valid( NastiArbiter_2_io_slave_aw_valid ),
       .io_slave_aw_bits_addr( NastiArbiter_2_io_slave_aw_bits_addr ),
       .io_slave_aw_bits_len( NastiArbiter_2_io_slave_aw_bits_len ),
       .io_slave_aw_bits_size( NastiArbiter_2_io_slave_aw_bits_size ),
       .io_slave_aw_bits_burst( NastiArbiter_2_io_slave_aw_bits_burst ),
       .io_slave_aw_bits_lock( NastiArbiter_2_io_slave_aw_bits_lock ),
       .io_slave_aw_bits_cache( NastiArbiter_2_io_slave_aw_bits_cache ),
       .io_slave_aw_bits_prot( NastiArbiter_2_io_slave_aw_bits_prot ),
       .io_slave_aw_bits_qos( NastiArbiter_2_io_slave_aw_bits_qos ),
       .io_slave_aw_bits_region( NastiArbiter_2_io_slave_aw_bits_region ),
       .io_slave_aw_bits_id( NastiArbiter_2_io_slave_aw_bits_id ),
       .io_slave_aw_bits_user( NastiArbiter_2_io_slave_aw_bits_user ),
       .io_slave_w_ready( io_slaves_2_w_ready ),
       .io_slave_w_valid( NastiArbiter_2_io_slave_w_valid ),
       .io_slave_w_bits_data( NastiArbiter_2_io_slave_w_bits_data ),
       .io_slave_w_bits_last( NastiArbiter_2_io_slave_w_bits_last ),
       .io_slave_w_bits_strb( NastiArbiter_2_io_slave_w_bits_strb ),
       .io_slave_w_bits_user( NastiArbiter_2_io_slave_w_bits_user ),
       .io_slave_b_ready( NastiArbiter_2_io_slave_b_ready ),
       .io_slave_b_valid( io_slaves_2_b_valid ),
       .io_slave_b_bits_resp( io_slaves_2_b_bits_resp ),
       .io_slave_b_bits_id( io_slaves_2_b_bits_id ),
       .io_slave_b_bits_user( io_slaves_2_b_bits_user ),
       .io_slave_ar_ready( io_slaves_2_ar_ready ),
       .io_slave_ar_valid( NastiArbiter_2_io_slave_ar_valid ),
       .io_slave_ar_bits_addr( NastiArbiter_2_io_slave_ar_bits_addr ),
       .io_slave_ar_bits_len( NastiArbiter_2_io_slave_ar_bits_len ),
       .io_slave_ar_bits_size( NastiArbiter_2_io_slave_ar_bits_size ),
       .io_slave_ar_bits_burst( NastiArbiter_2_io_slave_ar_bits_burst ),
       .io_slave_ar_bits_lock( NastiArbiter_2_io_slave_ar_bits_lock ),
       .io_slave_ar_bits_cache( NastiArbiter_2_io_slave_ar_bits_cache ),
       .io_slave_ar_bits_prot( NastiArbiter_2_io_slave_ar_bits_prot ),
       .io_slave_ar_bits_qos( NastiArbiter_2_io_slave_ar_bits_qos ),
       .io_slave_ar_bits_region( NastiArbiter_2_io_slave_ar_bits_region ),
       .io_slave_ar_bits_id( NastiArbiter_2_io_slave_ar_bits_id ),
       .io_slave_ar_bits_user( NastiArbiter_2_io_slave_ar_bits_user ),
       .io_slave_r_ready( NastiArbiter_2_io_slave_r_ready ),
       .io_slave_r_valid( io_slaves_2_r_valid ),
       .io_slave_r_bits_resp( io_slaves_2_r_bits_resp ),
       .io_slave_r_bits_data( io_slaves_2_r_bits_data ),
       .io_slave_r_bits_last( io_slaves_2_r_bits_last ),
       .io_slave_r_bits_id( io_slaves_2_r_bits_id ),
       .io_slave_r_bits_user( io_slaves_2_r_bits_user )
  );
endmodule

module NastiMultiChannelRouter(
    output io_master_aw_ready,
    input  io_master_aw_valid,
    input [31:0] io_master_aw_bits_addr,
    input [7:0] io_master_aw_bits_len,
    input [2:0] io_master_aw_bits_size,
    input [1:0] io_master_aw_bits_burst,
    input  io_master_aw_bits_lock,
    input [3:0] io_master_aw_bits_cache,
    input [2:0] io_master_aw_bits_prot,
    input [3:0] io_master_aw_bits_qos,
    input [3:0] io_master_aw_bits_region,
    input [4:0] io_master_aw_bits_id,
    input  io_master_aw_bits_user,
    output io_master_w_ready,
    input  io_master_w_valid,
    input [63:0] io_master_w_bits_data,
    input  io_master_w_bits_last,
    input [7:0] io_master_w_bits_strb,
    input  io_master_w_bits_user,
    input  io_master_b_ready,
    output io_master_b_valid,
    output[1:0] io_master_b_bits_resp,
    output[4:0] io_master_b_bits_id,
    output io_master_b_bits_user,
    output io_master_ar_ready,
    input  io_master_ar_valid,
    input [31:0] io_master_ar_bits_addr,
    input [7:0] io_master_ar_bits_len,
    input [2:0] io_master_ar_bits_size,
    input [1:0] io_master_ar_bits_burst,
    input  io_master_ar_bits_lock,
    input [3:0] io_master_ar_bits_cache,
    input [2:0] io_master_ar_bits_prot,
    input [3:0] io_master_ar_bits_qos,
    input [3:0] io_master_ar_bits_region,
    input [4:0] io_master_ar_bits_id,
    input  io_master_ar_bits_user,
    input  io_master_r_ready,
    output io_master_r_valid,
    output[1:0] io_master_r_bits_resp,
    output[63:0] io_master_r_bits_data,
    output io_master_r_bits_last,
    output[4:0] io_master_r_bits_id,
    output io_master_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[4:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [4:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[4:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [4:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);



  assign io_slaves_0_r_ready = io_master_r_ready;
  assign io_slaves_0_ar_bits_user = io_master_ar_bits_user;
  assign io_slaves_0_ar_bits_id = io_master_ar_bits_id;
  assign io_slaves_0_ar_bits_region = io_master_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = io_master_ar_bits_size;
  assign io_slaves_0_ar_bits_len = io_master_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slaves_0_ar_valid = io_master_ar_valid;
  assign io_slaves_0_b_ready = io_master_b_ready;
  assign io_slaves_0_w_bits_user = io_master_w_bits_user;
  assign io_slaves_0_w_bits_strb = io_master_w_bits_strb;
  assign io_slaves_0_w_bits_last = io_master_w_bits_last;
  assign io_slaves_0_w_bits_data = io_master_w_bits_data;
  assign io_slaves_0_w_valid = io_master_w_valid;
  assign io_slaves_0_aw_bits_user = io_master_aw_bits_user;
  assign io_slaves_0_aw_bits_id = io_master_aw_bits_id;
  assign io_slaves_0_aw_bits_region = io_master_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = io_master_aw_bits_size;
  assign io_slaves_0_aw_bits_len = io_master_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slaves_0_aw_valid = io_master_aw_valid;
  assign io_master_r_bits_user = io_slaves_0_r_bits_user;
  assign io_master_r_bits_id = io_slaves_0_r_bits_id;
  assign io_master_r_bits_last = io_slaves_0_r_bits_last;
  assign io_master_r_bits_data = io_slaves_0_r_bits_data;
  assign io_master_r_bits_resp = io_slaves_0_r_bits_resp;
  assign io_master_r_valid = io_slaves_0_r_valid;
  assign io_master_ar_ready = io_slaves_0_ar_ready;
  assign io_master_b_bits_user = io_slaves_0_b_bits_user;
  assign io_master_b_bits_id = io_slaves_0_b_bits_id;
  assign io_master_b_bits_resp = io_slaves_0_b_bits_resp;
  assign io_master_b_valid = io_slaves_0_b_valid;
  assign io_master_w_ready = io_slaves_0_w_ready;
  assign io_master_aw_ready = io_slaves_0_aw_ready;
endmodule

module RRArbiter_6(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [4:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [4:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [4:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[4:0] io_out_bits_id,
    output io_out_bits_user,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire T3;
  wire T4;
  reg [1:0] last_grant;
  wire[1:0] T58;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[1:0] T12;
  wire T13;
  wire[4:0] T14;
  wire[4:0] T15;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T7 ? 2'h1 : T0;
  assign T0 = T3 ? 2'h2 : T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T3 = io_in_2_valid & T4;
  assign T4 = last_grant < 2'h2;
  assign T58 = reset ? 2'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = io_in_1_valid & T8;
  assign T8 = last_grant < 2'h1;
  assign io_out_bits_user = T9;
  assign T9 = T13 ? io_in_2_bits_user : T10;
  assign T10 = T11 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = chosen;
  assign T13 = T12[1'h1:1'h1];
  assign io_out_bits_id = T14;
  assign T14 = T17 ? io_in_2_bits_id : T15;
  assign T15 = T16 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T16 = T12[1'h0:1'h0];
  assign T17 = T12[1'h1:1'h1];
  assign io_out_bits_resp = T18;
  assign T18 = T21 ? io_in_2_bits_resp : T19;
  assign T19 = T20 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign io_out_valid = T22;
  assign T22 = T25 ? io_in_2_valid : T23;
  assign T23 = T24 ? io_in_1_valid : io_in_0_valid;
  assign T24 = T12[1'h0:1'h0];
  assign T25 = T12[1'h1:1'h1];
  assign io_in_0_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T37 | T28;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T32 | T30;
  assign T30 = io_in_2_valid & T31;
  assign T31 = last_grant < 2'h2;
  assign T32 = T35 | T33;
  assign T33 = io_in_1_valid & T34;
  assign T34 = last_grant < 2'h1;
  assign T35 = io_in_0_valid & T36;
  assign T36 = last_grant < 2'h0;
  assign T37 = last_grant < 2'h0;
  assign io_in_1_ready = T38;
  assign T38 = T39 & io_out_ready;
  assign T39 = T44 | T40;
  assign T40 = T41 ^ 1'h1;
  assign T41 = T42 | io_in_0_valid;
  assign T42 = T43 | T30;
  assign T43 = T35 | T33;
  assign T44 = T46 & T45;
  assign T45 = last_grant < 2'h1;
  assign T46 = T35 ^ 1'h1;
  assign io_in_2_ready = T47;
  assign T47 = T48 & io_out_ready;
  assign T48 = T54 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_1_valid;
  assign T51 = T52 | io_in_0_valid;
  assign T52 = T53 | T30;
  assign T53 = T35 | T33;
  assign T54 = T56 & T55;
  assign T55 = last_grant < 2'h2;
  assign T56 = T57 ^ 1'h1;
  assign T57 = T35 | T33;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module JunctionsPeekingArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [63:0] io_in_2_bits_data,
    input  io_in_2_bits_last,
    input [4:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [63:0] io_in_1_bits_data,
    input  io_in_1_bits_last,
    input [4:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_last,
    input [4:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[63:0] io_out_bits_data,
    output io_out_bits_last,
    output[4:0] io_out_bits_id,
    output io_out_bits_user
);

  wire T0;
  wire T1;
  wire T2;
  wire[1:0] T3;
  wire[1:0] chosen;
  wire[1:0] choice;
  wire[1:0] T4;
  wire[1:0] T5;
  reg [1:0] T6;
  wire[1:0] T8;
  wire[1:0] T9;
  reg [1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire[1:0] T13;
  reg [1:0] T14;
  wire[1:0] T15;
  reg [1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire[1:0] T34;
  reg [1:0] T35;
  wire[1:0] T36;
  reg [1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  reg [1:0] lockIdx;
  wire[1:0] T88;
  wire[1:0] T54;
  wire T55;
  wire T56;
  wire T57;
  reg  locked;
  wire T89;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[4:0] T62;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[63:0] T70;
  wire[63:0] T71;
  wire T72;
  wire T73;
  wire[1:0] T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_bits_user = T0;
  assign T0 = T61 ? io_in_2_bits_user : T1;
  assign T1 = T2 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T2 = T3[1'h0:1'h0];
  assign T3 = chosen;
  assign chosen = locked ? lockIdx : choice;
  assign choice = T40 ? T34 : T4;
  assign T4 = T19 ? T13 : T5;
  assign T5 = T12 ? T10 : T6;
  always @(*) case (T8)
    0: T6 = 2'h0;
    1: T6 = 2'h1;
    2: T6 = 2'h2;
    default: begin
      T6 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T6 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T8 = T9 - 2'h1;
  assign T9 = lockIdx + 2'h1;
  always @(*) case (T11)
    0: T10 = 2'h0;
    1: T10 = 2'h1;
    2: T10 = 2'h2;
    default: begin
      T10 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T10 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T11 = 2'h2 + T9;
  assign T12 = T9 < 2'h1;
  assign T13 = T18 ? T16 : T14;
  always @(*) case (T15)
    0: T14 = 2'h0;
    1: T14 = 2'h1;
    2: T14 = 2'h2;
    default: begin
      T14 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T14 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T15 = T9 - 2'h2;
  always @(*) case (T17)
    0: T16 = 2'h0;
    1: T16 = 2'h1;
    2: T16 = 2'h2;
    default: begin
      T16 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T16 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T17 = 2'h1 + T9;
  assign T18 = T9 < 2'h2;
  assign T19 = T33 ? T27 : T20;
  assign T20 = T26 ? io_in_2_valid : T21;
  assign T21 = T22 ? io_in_1_valid : io_in_0_valid;
  assign T22 = T23[1'h0:1'h0];
  assign T23 = T24;
  assign T24 = T25 - 2'h2;
  assign T25 = lockIdx + 2'h1;
  assign T26 = T23[1'h1:1'h1];
  assign T27 = T32 ? io_in_2_valid : T28;
  assign T28 = T29 ? io_in_1_valid : io_in_0_valid;
  assign T29 = T30[1'h0:1'h0];
  assign T30 = T31;
  assign T31 = 2'h1 + T25;
  assign T32 = T30[1'h1:1'h1];
  assign T33 = T25 < 2'h2;
  assign T34 = T39 ? T37 : T35;
  always @(*) case (T36)
    0: T35 = 2'h0;
    1: T35 = 2'h1;
    2: T35 = 2'h2;
    default: begin
      T35 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T35 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T36 = T9 - 2'h3;
  always @(*) case (T38)
    0: T37 = 2'h0;
    1: T37 = 2'h1;
    2: T37 = 2'h2;
    default: begin
      T37 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T37 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T38 = 2'h0 + T9;
  assign T39 = T9 < 2'h3;
  assign T40 = T53 ? T47 : T41;
  assign T41 = T46 ? io_in_2_valid : T42;
  assign T42 = T43 ? io_in_1_valid : io_in_0_valid;
  assign T43 = T44[1'h0:1'h0];
  assign T44 = T45;
  assign T45 = T25 - 2'h3;
  assign T46 = T44[1'h1:1'h1];
  assign T47 = T52 ? io_in_2_valid : T48;
  assign T48 = T49 ? io_in_1_valid : io_in_0_valid;
  assign T49 = T50[1'h0:1'h0];
  assign T50 = T51;
  assign T51 = 2'h0 + T25;
  assign T52 = T50[1'h1:1'h1];
  assign T53 = T25 < 2'h3;
  assign T88 = reset ? 2'h0 : T54;
  assign T54 = T55 ? choice : lockIdx;
  assign T55 = T57 & T56;
  assign T56 = locked ^ 1'h1;
  assign T57 = io_out_ready & io_out_valid;
  assign T89 = reset ? 1'h0 : T58;
  assign T58 = T60 ? 1'h0 : T59;
  assign T59 = T55 ? 1'h1 : locked;
  assign T60 = T57 & io_out_bits_last;
  assign T61 = T3[1'h1:1'h1];
  assign io_out_bits_id = T62;
  assign T62 = T65 ? io_in_2_bits_id : T63;
  assign T63 = T64 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T64 = T3[1'h0:1'h0];
  assign T65 = T3[1'h1:1'h1];
  assign io_out_bits_last = T66;
  assign T66 = T69 ? io_in_2_bits_last : T67;
  assign T67 = T68 ? io_in_1_bits_last : io_in_0_bits_last;
  assign T68 = T3[1'h0:1'h0];
  assign T69 = T3[1'h1:1'h1];
  assign io_out_bits_data = T70;
  assign T70 = T73 ? io_in_2_bits_data : T71;
  assign T71 = T72 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T72 = T3[1'h0:1'h0];
  assign T73 = T3[1'h1:1'h1];
  assign io_out_bits_resp = T74;
  assign T74 = T77 ? io_in_2_bits_resp : T75;
  assign T75 = T76 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T76 = T3[1'h0:1'h0];
  assign T77 = T3[1'h1:1'h1];
  assign io_out_valid = T78;
  assign T78 = T81 ? io_in_2_valid : T79;
  assign T79 = T80 ? io_in_1_valid : io_in_0_valid;
  assign T80 = T3[1'h0:1'h0];
  assign T81 = T3[1'h1:1'h1];
  assign io_in_0_ready = T82;
  assign T82 = io_out_ready & T83;
  assign T83 = chosen == 2'h0;
  assign io_in_1_ready = T84;
  assign T84 = io_out_ready & T85;
  assign T85 = chosen == 2'h1;
  assign io_in_2_ready = T86;
  assign T86 = io_out_ready & T87;
  assign T87 = chosen == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 2'h0;
    end else if(T55) begin
      lockIdx <= choice;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T60) begin
      locked <= 1'h0;
    end else if(T55) begin
      locked <= 1'h1;
    end
  end
endmodule

module NastiRouter_1(input clk, input reset,
    output io_master_aw_ready,
    input  io_master_aw_valid,
    input [31:0] io_master_aw_bits_addr,
    input [7:0] io_master_aw_bits_len,
    input [2:0] io_master_aw_bits_size,
    input [1:0] io_master_aw_bits_burst,
    input  io_master_aw_bits_lock,
    input [3:0] io_master_aw_bits_cache,
    input [2:0] io_master_aw_bits_prot,
    input [3:0] io_master_aw_bits_qos,
    input [3:0] io_master_aw_bits_region,
    input [4:0] io_master_aw_bits_id,
    input  io_master_aw_bits_user,
    output io_master_w_ready,
    input  io_master_w_valid,
    input [63:0] io_master_w_bits_data,
    input  io_master_w_bits_last,
    input [7:0] io_master_w_bits_strb,
    input  io_master_w_bits_user,
    input  io_master_b_ready,
    output io_master_b_valid,
    output[1:0] io_master_b_bits_resp,
    output[4:0] io_master_b_bits_id,
    output io_master_b_bits_user,
    output io_master_ar_ready,
    input  io_master_ar_valid,
    input [31:0] io_master_ar_bits_addr,
    input [7:0] io_master_ar_bits_len,
    input [2:0] io_master_ar_bits_size,
    input [1:0] io_master_ar_bits_burst,
    input  io_master_ar_bits_lock,
    input [3:0] io_master_ar_bits_cache,
    input [2:0] io_master_ar_bits_prot,
    input [3:0] io_master_ar_bits_qos,
    input [3:0] io_master_ar_bits_region,
    input [4:0] io_master_ar_bits_id,
    input  io_master_ar_bits_user,
    input  io_master_r_ready,
    output io_master_r_valid,
    output[1:0] io_master_r_bits_resp,
    output[63:0] io_master_r_bits_data,
    output io_master_r_bits_last,
    output[4:0] io_master_r_bits_id,
    output io_master_r_bits_user,
    input  io_slave_1_aw_ready,
    output io_slave_1_aw_valid,
    output[31:0] io_slave_1_aw_bits_addr,
    output[7:0] io_slave_1_aw_bits_len,
    output[2:0] io_slave_1_aw_bits_size,
    output[1:0] io_slave_1_aw_bits_burst,
    output io_slave_1_aw_bits_lock,
    output[3:0] io_slave_1_aw_bits_cache,
    output[2:0] io_slave_1_aw_bits_prot,
    output[3:0] io_slave_1_aw_bits_qos,
    output[3:0] io_slave_1_aw_bits_region,
    output[4:0] io_slave_1_aw_bits_id,
    output io_slave_1_aw_bits_user,
    input  io_slave_1_w_ready,
    output io_slave_1_w_valid,
    output[63:0] io_slave_1_w_bits_data,
    output io_slave_1_w_bits_last,
    output[7:0] io_slave_1_w_bits_strb,
    output io_slave_1_w_bits_user,
    output io_slave_1_b_ready,
    input  io_slave_1_b_valid,
    input [1:0] io_slave_1_b_bits_resp,
    input [4:0] io_slave_1_b_bits_id,
    input  io_slave_1_b_bits_user,
    input  io_slave_1_ar_ready,
    output io_slave_1_ar_valid,
    output[31:0] io_slave_1_ar_bits_addr,
    output[7:0] io_slave_1_ar_bits_len,
    output[2:0] io_slave_1_ar_bits_size,
    output[1:0] io_slave_1_ar_bits_burst,
    output io_slave_1_ar_bits_lock,
    output[3:0] io_slave_1_ar_bits_cache,
    output[2:0] io_slave_1_ar_bits_prot,
    output[3:0] io_slave_1_ar_bits_qos,
    output[3:0] io_slave_1_ar_bits_region,
    output[4:0] io_slave_1_ar_bits_id,
    output io_slave_1_ar_bits_user,
    output io_slave_1_r_ready,
    input  io_slave_1_r_valid,
    input [1:0] io_slave_1_r_bits_resp,
    input [63:0] io_slave_1_r_bits_data,
    input  io_slave_1_r_bits_last,
    input [4:0] io_slave_1_r_bits_id,
    input  io_slave_1_r_bits_user,
    input  io_slave_0_aw_ready,
    output io_slave_0_aw_valid,
    output[31:0] io_slave_0_aw_bits_addr,
    output[7:0] io_slave_0_aw_bits_len,
    output[2:0] io_slave_0_aw_bits_size,
    output[1:0] io_slave_0_aw_bits_burst,
    output io_slave_0_aw_bits_lock,
    output[3:0] io_slave_0_aw_bits_cache,
    output[2:0] io_slave_0_aw_bits_prot,
    output[3:0] io_slave_0_aw_bits_qos,
    output[3:0] io_slave_0_aw_bits_region,
    output[4:0] io_slave_0_aw_bits_id,
    output io_slave_0_aw_bits_user,
    input  io_slave_0_w_ready,
    output io_slave_0_w_valid,
    output[63:0] io_slave_0_w_bits_data,
    output io_slave_0_w_bits_last,
    output[7:0] io_slave_0_w_bits_strb,
    output io_slave_0_w_bits_user,
    output io_slave_0_b_ready,
    input  io_slave_0_b_valid,
    input [1:0] io_slave_0_b_bits_resp,
    input [4:0] io_slave_0_b_bits_id,
    input  io_slave_0_b_bits_user,
    input  io_slave_0_ar_ready,
    output io_slave_0_ar_valid,
    output[31:0] io_slave_0_ar_bits_addr,
    output[7:0] io_slave_0_ar_bits_len,
    output[2:0] io_slave_0_ar_bits_size,
    output[1:0] io_slave_0_ar_bits_burst,
    output io_slave_0_ar_bits_lock,
    output[3:0] io_slave_0_ar_bits_cache,
    output[2:0] io_slave_0_ar_bits_prot,
    output[3:0] io_slave_0_ar_bits_qos,
    output[3:0] io_slave_0_ar_bits_region,
    output[4:0] io_slave_0_ar_bits_id,
    output io_slave_0_ar_bits_user,
    output io_slave_0_r_ready,
    input  io_slave_0_r_valid,
    input [1:0] io_slave_0_r_bits_resp,
    input [63:0] io_slave_0_r_bits_data,
    input  io_slave_0_r_bits_last,
    input [4:0] io_slave_0_r_bits_id,
    input  io_slave_0_r_bits_user
);

  wire T0;
  wire r_invalid;
  wire T1;
  wire[1:0] ar_route;
  wire[1:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire w_invalid;
  wire T10;
  wire[1:0] aw_route;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg  R21;
  wire T55;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  R32;
  wire T56;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire ar_ready;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire w_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire aw_ready;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire b_arb_io_in_2_ready;
  wire b_arb_io_in_1_ready;
  wire b_arb_io_in_0_ready;
  wire b_arb_io_out_valid;
  wire[1:0] b_arb_io_out_bits_resp;
  wire[4:0] b_arb_io_out_bits_id;
  wire b_arb_io_out_bits_user;
  wire r_arb_io_in_2_ready;
  wire r_arb_io_in_1_ready;
  wire r_arb_io_in_0_ready;
  wire r_arb_io_out_valid;
  wire[1:0] r_arb_io_out_bits_resp;
  wire[63:0] r_arb_io_out_bits_data;
  wire r_arb_io_out_bits_last;
  wire[4:0] r_arb_io_out_bits_id;
  wire r_arb_io_out_bits_user;
  wire err_slave_io_aw_ready;
  wire err_slave_io_w_ready;
  wire err_slave_io_b_valid;
  wire[1:0] err_slave_io_b_bits_resp;
  wire[4:0] err_slave_io_b_bits_id;
  wire err_slave_io_ar_ready;
  wire err_slave_io_r_valid;
  wire[1:0] err_slave_io_r_bits_resp;
  wire[63:0] err_slave_io_r_bits_data;
  wire err_slave_io_r_bits_last;
  wire[4:0] err_slave_io_r_bits_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R21 = {1{$random}};
    R32 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = r_invalid & io_master_ar_valid;
  assign r_invalid = T1 ^ 1'h1;
  assign T1 = ar_route != 2'h0;
  assign ar_route = T2;
  assign T2 = {T6, T3};
  assign T3 = T5 & T4;
  assign T4 = io_master_ar_bits_addr < 32'h40008000;
  assign T5 = 32'h40000000 <= io_master_ar_bits_addr;
  assign T6 = T8 & T7;
  assign T7 = io_master_ar_bits_addr < 32'h40008200;
  assign T8 = 32'h40008000 <= io_master_ar_bits_addr;
  assign T9 = w_invalid & io_master_aw_valid;
  assign w_invalid = T10 ^ 1'h1;
  assign T10 = aw_route != 2'h0;
  assign aw_route = T11;
  assign T11 = {T15, T12};
  assign T12 = T14 & T13;
  assign T13 = io_master_aw_bits_addr < 32'h40008000;
  assign T14 = 32'h40000000 <= io_master_aw_bits_addr;
  assign T15 = T17 & T16;
  assign T16 = io_master_aw_bits_addr < 32'h40008200;
  assign T17 = 32'h40008000 <= io_master_aw_bits_addr;
  assign io_slave_0_r_ready = r_arb_io_in_0_ready;
  assign io_slave_0_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_0_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_0_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_0_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_0_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_0_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_0_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_0_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_0_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_0_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_0_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_0_ar_valid = T18;
  assign T18 = io_master_ar_valid & T19;
  assign T19 = ar_route[1'h0:1'h0];
  assign io_slave_0_b_ready = b_arb_io_in_0_ready;
  assign io_slave_0_w_bits_user = io_master_w_bits_user;
  assign io_slave_0_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_0_w_bits_last = io_master_w_bits_last;
  assign io_slave_0_w_bits_data = io_master_w_bits_data;
  assign io_slave_0_w_valid = T20;
  assign T20 = io_master_w_valid & R21;
  assign T55 = reset ? 1'h0 : T22;
  assign T22 = T25 ? 1'h0 : T23;
  assign T23 = T24 ? 1'h1 : R21;
  assign T24 = io_slave_0_aw_ready & io_slave_0_aw_valid;
  assign T25 = T26 & io_slave_0_w_bits_last;
  assign T26 = io_slave_0_w_ready & io_slave_0_w_valid;
  assign io_slave_0_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_0_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_0_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_0_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_0_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_0_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_0_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_0_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_0_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_0_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_0_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_0_aw_valid = T27;
  assign T27 = io_master_aw_valid & T28;
  assign T28 = aw_route[1'h0:1'h0];
  assign io_slave_1_r_ready = r_arb_io_in_1_ready;
  assign io_slave_1_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_1_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_1_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_1_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_1_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_1_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_1_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_1_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_1_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_1_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_1_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_1_ar_valid = T29;
  assign T29 = io_master_ar_valid & T30;
  assign T30 = ar_route[1'h1:1'h1];
  assign io_slave_1_b_ready = b_arb_io_in_1_ready;
  assign io_slave_1_w_bits_user = io_master_w_bits_user;
  assign io_slave_1_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_1_w_bits_last = io_master_w_bits_last;
  assign io_slave_1_w_bits_data = io_master_w_bits_data;
  assign io_slave_1_w_valid = T31;
  assign T31 = io_master_w_valid & R32;
  assign T56 = reset ? 1'h0 : T33;
  assign T33 = T36 ? 1'h0 : T34;
  assign T34 = T35 ? 1'h1 : R32;
  assign T35 = io_slave_1_aw_ready & io_slave_1_aw_valid;
  assign T36 = T37 & io_slave_1_w_bits_last;
  assign T37 = io_slave_1_w_ready & io_slave_1_w_valid;
  assign io_slave_1_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_1_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_1_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_1_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_1_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_1_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_1_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_1_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_1_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_1_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_1_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_1_aw_valid = T38;
  assign T38 = io_master_aw_valid & T39;
  assign T39 = aw_route[1'h1:1'h1];
  assign io_master_r_bits_user = r_arb_io_out_bits_user;
  assign io_master_r_bits_id = r_arb_io_out_bits_id;
  assign io_master_r_bits_last = r_arb_io_out_bits_last;
  assign io_master_r_bits_data = r_arb_io_out_bits_data;
  assign io_master_r_bits_resp = r_arb_io_out_bits_resp;
  assign io_master_r_valid = r_arb_io_out_valid;
  assign io_master_ar_ready = T40;
  assign T40 = ar_ready | T41;
  assign T41 = r_invalid & err_slave_io_ar_ready;
  assign ar_ready = T44 | T42;
  assign T42 = io_slave_1_ar_ready & T43;
  assign T43 = ar_route[1'h1:1'h1];
  assign T44 = io_slave_0_ar_ready & T45;
  assign T45 = ar_route[1'h0:1'h0];
  assign io_master_b_bits_user = b_arb_io_out_bits_user;
  assign io_master_b_bits_id = b_arb_io_out_bits_id;
  assign io_master_b_bits_resp = b_arb_io_out_bits_resp;
  assign io_master_b_valid = b_arb_io_out_valid;
  assign io_master_w_ready = T46;
  assign T46 = w_ready | err_slave_io_w_ready;
  assign w_ready = T48 | T47;
  assign T47 = io_slave_1_w_ready & R32;
  assign T48 = io_slave_0_w_ready & R21;
  assign io_master_aw_ready = T49;
  assign T49 = aw_ready | T50;
  assign T50 = w_invalid & err_slave_io_aw_ready;
  assign aw_ready = T53 | T51;
  assign T51 = io_slave_1_aw_ready & T52;
  assign T52 = aw_route[1'h1:1'h1];
  assign T53 = io_slave_0_aw_ready & T54;
  assign T54 = aw_route[1'h0:1'h0];
  NastiErrorSlave err_slave(.clk(clk), .reset(reset),
       .io_aw_ready( err_slave_io_aw_ready ),
       .io_aw_valid( T9 ),
       .io_aw_bits_addr( io_master_aw_bits_addr ),
       .io_aw_bits_len( io_master_aw_bits_len ),
       .io_aw_bits_size( io_master_aw_bits_size ),
       .io_aw_bits_burst( io_master_aw_bits_burst ),
       .io_aw_bits_lock( io_master_aw_bits_lock ),
       .io_aw_bits_cache( io_master_aw_bits_cache ),
       .io_aw_bits_prot( io_master_aw_bits_prot ),
       .io_aw_bits_qos( io_master_aw_bits_qos ),
       .io_aw_bits_region( io_master_aw_bits_region ),
       .io_aw_bits_id( io_master_aw_bits_id ),
       .io_aw_bits_user( io_master_aw_bits_user ),
       .io_w_ready( err_slave_io_w_ready ),
       .io_w_valid( io_master_w_valid ),
       .io_w_bits_data( io_master_w_bits_data ),
       .io_w_bits_last( io_master_w_bits_last ),
       .io_w_bits_strb( io_master_w_bits_strb ),
       .io_w_bits_user( io_master_w_bits_user ),
       .io_b_ready( b_arb_io_in_2_ready ),
       .io_b_valid( err_slave_io_b_valid ),
       .io_b_bits_resp( err_slave_io_b_bits_resp ),
       .io_b_bits_id( err_slave_io_b_bits_id ),
       //.io_b_bits_user(  )
       .io_ar_ready( err_slave_io_ar_ready ),
       .io_ar_valid( T0 ),
       .io_ar_bits_addr( io_master_ar_bits_addr ),
       .io_ar_bits_len( io_master_ar_bits_len ),
       .io_ar_bits_size( io_master_ar_bits_size ),
       .io_ar_bits_burst( io_master_ar_bits_burst ),
       .io_ar_bits_lock( io_master_ar_bits_lock ),
       .io_ar_bits_cache( io_master_ar_bits_cache ),
       .io_ar_bits_prot( io_master_ar_bits_prot ),
       .io_ar_bits_qos( io_master_ar_bits_qos ),
       .io_ar_bits_region( io_master_ar_bits_region ),
       .io_ar_bits_id( io_master_ar_bits_id ),
       .io_ar_bits_user( io_master_ar_bits_user ),
       .io_r_ready( r_arb_io_in_2_ready ),
       .io_r_valid( err_slave_io_r_valid ),
       .io_r_bits_resp( err_slave_io_r_bits_resp ),
       .io_r_bits_data( err_slave_io_r_bits_data ),
       .io_r_bits_last( err_slave_io_r_bits_last ),
       .io_r_bits_id( err_slave_io_r_bits_id )
       //.io_r_bits_user(  )
  );
  RRArbiter_6 b_arb(.clk(clk), .reset(reset),
       .io_in_2_ready( b_arb_io_in_2_ready ),
       .io_in_2_valid( err_slave_io_b_valid ),
       .io_in_2_bits_resp( err_slave_io_b_bits_resp ),
       .io_in_2_bits_id( err_slave_io_b_bits_id ),
       //.io_in_2_bits_user(  )
       .io_in_1_ready( b_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_b_valid ),
       .io_in_1_bits_resp( io_slave_1_b_bits_resp ),
       .io_in_1_bits_id( io_slave_1_b_bits_id ),
       .io_in_1_bits_user( io_slave_1_b_bits_user ),
       .io_in_0_ready( b_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_b_valid ),
       .io_in_0_bits_resp( io_slave_0_b_bits_resp ),
       .io_in_0_bits_id( io_slave_0_b_bits_id ),
       .io_in_0_bits_user( io_slave_0_b_bits_user ),
       .io_out_ready( io_master_b_ready ),
       .io_out_valid( b_arb_io_out_valid ),
       .io_out_bits_resp( b_arb_io_out_bits_resp ),
       .io_out_bits_id( b_arb_io_out_bits_id ),
       .io_out_bits_user( b_arb_io_out_bits_user )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign b_arb.io_in_2_bits_user = {1{$random}};
// synthesis translate_on
`endif
  JunctionsPeekingArbiter_1 r_arb(.clk(clk), .reset(reset),
       .io_in_2_ready( r_arb_io_in_2_ready ),
       .io_in_2_valid( err_slave_io_r_valid ),
       .io_in_2_bits_resp( err_slave_io_r_bits_resp ),
       .io_in_2_bits_data( err_slave_io_r_bits_data ),
       .io_in_2_bits_last( err_slave_io_r_bits_last ),
       .io_in_2_bits_id( err_slave_io_r_bits_id ),
       //.io_in_2_bits_user(  )
       .io_in_1_ready( r_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_r_valid ),
       .io_in_1_bits_resp( io_slave_1_r_bits_resp ),
       .io_in_1_bits_data( io_slave_1_r_bits_data ),
       .io_in_1_bits_last( io_slave_1_r_bits_last ),
       .io_in_1_bits_id( io_slave_1_r_bits_id ),
       .io_in_1_bits_user( io_slave_1_r_bits_user ),
       .io_in_0_ready( r_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_r_valid ),
       .io_in_0_bits_resp( io_slave_0_r_bits_resp ),
       .io_in_0_bits_data( io_slave_0_r_bits_data ),
       .io_in_0_bits_last( io_slave_0_r_bits_last ),
       .io_in_0_bits_id( io_slave_0_r_bits_id ),
       .io_in_0_bits_user( io_slave_0_r_bits_user ),
       .io_out_ready( io_master_r_ready ),
       .io_out_valid( r_arb_io_out_valid ),
       .io_out_bits_resp( r_arb_io_out_bits_resp ),
       .io_out_bits_data( r_arb_io_out_bits_data ),
       .io_out_bits_last( r_arb_io_out_bits_last ),
       .io_out_bits_id( r_arb_io_out_bits_id ),
       .io_out_bits_user( r_arb_io_out_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign r_arb.io_in_2_bits_user = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      R21 <= 1'h0;
    end else if(T25) begin
      R21 <= 1'h0;
    end else if(T24) begin
      R21 <= 1'h1;
    end
    if(reset) begin
      R32 <= 1'h0;
    end else if(T36) begin
      R32 <= 1'h0;
    end else if(T35) begin
      R32 <= 1'h1;
    end
  end
endmodule

module NastiCrossbar_1(input clk, input reset,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [4:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[4:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [4:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[4:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[4:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [4:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[4:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [4:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[4:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [4:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[4:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [4:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire NastiRouter_io_master_aw_ready;
  wire NastiRouter_io_master_w_ready;
  wire NastiRouter_io_master_b_valid;
  wire[1:0] NastiRouter_io_master_b_bits_resp;
  wire[4:0] NastiRouter_io_master_b_bits_id;
  wire NastiRouter_io_master_b_bits_user;
  wire NastiRouter_io_master_ar_ready;
  wire NastiRouter_io_master_r_valid;
  wire[1:0] NastiRouter_io_master_r_bits_resp;
  wire[63:0] NastiRouter_io_master_r_bits_data;
  wire NastiRouter_io_master_r_bits_last;
  wire[4:0] NastiRouter_io_master_r_bits_id;
  wire NastiRouter_io_master_r_bits_user;
  wire NastiRouter_io_slave_1_aw_valid;
  wire[31:0] NastiRouter_io_slave_1_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_1_aw_bits_burst;
  wire NastiRouter_io_slave_1_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_region;
  wire[4:0] NastiRouter_io_slave_1_aw_bits_id;
  wire NastiRouter_io_slave_1_aw_bits_user;
  wire NastiRouter_io_slave_1_w_valid;
  wire[63:0] NastiRouter_io_slave_1_w_bits_data;
  wire NastiRouter_io_slave_1_w_bits_last;
  wire[7:0] NastiRouter_io_slave_1_w_bits_strb;
  wire NastiRouter_io_slave_1_w_bits_user;
  wire NastiRouter_io_slave_1_b_ready;
  wire NastiRouter_io_slave_1_ar_valid;
  wire[31:0] NastiRouter_io_slave_1_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_1_ar_bits_burst;
  wire NastiRouter_io_slave_1_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_region;
  wire[4:0] NastiRouter_io_slave_1_ar_bits_id;
  wire NastiRouter_io_slave_1_ar_bits_user;
  wire NastiRouter_io_slave_1_r_ready;
  wire NastiRouter_io_slave_0_aw_valid;
  wire[31:0] NastiRouter_io_slave_0_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_0_aw_bits_burst;
  wire NastiRouter_io_slave_0_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_region;
  wire[4:0] NastiRouter_io_slave_0_aw_bits_id;
  wire NastiRouter_io_slave_0_aw_bits_user;
  wire NastiRouter_io_slave_0_w_valid;
  wire[63:0] NastiRouter_io_slave_0_w_bits_data;
  wire NastiRouter_io_slave_0_w_bits_last;
  wire[7:0] NastiRouter_io_slave_0_w_bits_strb;
  wire NastiRouter_io_slave_0_w_bits_user;
  wire NastiRouter_io_slave_0_b_ready;
  wire NastiRouter_io_slave_0_ar_valid;
  wire[31:0] NastiRouter_io_slave_0_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_0_ar_bits_burst;
  wire NastiRouter_io_slave_0_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_region;
  wire[4:0] NastiRouter_io_slave_0_ar_bits_id;
  wire NastiRouter_io_slave_0_ar_bits_user;
  wire NastiRouter_io_slave_0_r_ready;


  assign io_slaves_0_r_ready = NastiRouter_io_slave_0_r_ready;
  assign io_slaves_0_ar_bits_user = NastiRouter_io_slave_0_ar_bits_user;
  assign io_slaves_0_ar_bits_id = NastiRouter_io_slave_0_ar_bits_id;
  assign io_slaves_0_ar_bits_region = NastiRouter_io_slave_0_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = NastiRouter_io_slave_0_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = NastiRouter_io_slave_0_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = NastiRouter_io_slave_0_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = NastiRouter_io_slave_0_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = NastiRouter_io_slave_0_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = NastiRouter_io_slave_0_ar_bits_size;
  assign io_slaves_0_ar_bits_len = NastiRouter_io_slave_0_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = NastiRouter_io_slave_0_ar_bits_addr;
  assign io_slaves_0_ar_valid = NastiRouter_io_slave_0_ar_valid;
  assign io_slaves_0_b_ready = NastiRouter_io_slave_0_b_ready;
  assign io_slaves_0_w_bits_user = NastiRouter_io_slave_0_w_bits_user;
  assign io_slaves_0_w_bits_strb = NastiRouter_io_slave_0_w_bits_strb;
  assign io_slaves_0_w_bits_last = NastiRouter_io_slave_0_w_bits_last;
  assign io_slaves_0_w_bits_data = NastiRouter_io_slave_0_w_bits_data;
  assign io_slaves_0_w_valid = NastiRouter_io_slave_0_w_valid;
  assign io_slaves_0_aw_bits_user = NastiRouter_io_slave_0_aw_bits_user;
  assign io_slaves_0_aw_bits_id = NastiRouter_io_slave_0_aw_bits_id;
  assign io_slaves_0_aw_bits_region = NastiRouter_io_slave_0_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = NastiRouter_io_slave_0_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = NastiRouter_io_slave_0_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = NastiRouter_io_slave_0_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = NastiRouter_io_slave_0_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = NastiRouter_io_slave_0_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = NastiRouter_io_slave_0_aw_bits_size;
  assign io_slaves_0_aw_bits_len = NastiRouter_io_slave_0_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = NastiRouter_io_slave_0_aw_bits_addr;
  assign io_slaves_0_aw_valid = NastiRouter_io_slave_0_aw_valid;
  assign io_slaves_1_r_ready = NastiRouter_io_slave_1_r_ready;
  assign io_slaves_1_ar_bits_user = NastiRouter_io_slave_1_ar_bits_user;
  assign io_slaves_1_ar_bits_id = NastiRouter_io_slave_1_ar_bits_id;
  assign io_slaves_1_ar_bits_region = NastiRouter_io_slave_1_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = NastiRouter_io_slave_1_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = NastiRouter_io_slave_1_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = NastiRouter_io_slave_1_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = NastiRouter_io_slave_1_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = NastiRouter_io_slave_1_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = NastiRouter_io_slave_1_ar_bits_size;
  assign io_slaves_1_ar_bits_len = NastiRouter_io_slave_1_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = NastiRouter_io_slave_1_ar_bits_addr;
  assign io_slaves_1_ar_valid = NastiRouter_io_slave_1_ar_valid;
  assign io_slaves_1_b_ready = NastiRouter_io_slave_1_b_ready;
  assign io_slaves_1_w_bits_user = NastiRouter_io_slave_1_w_bits_user;
  assign io_slaves_1_w_bits_strb = NastiRouter_io_slave_1_w_bits_strb;
  assign io_slaves_1_w_bits_last = NastiRouter_io_slave_1_w_bits_last;
  assign io_slaves_1_w_bits_data = NastiRouter_io_slave_1_w_bits_data;
  assign io_slaves_1_w_valid = NastiRouter_io_slave_1_w_valid;
  assign io_slaves_1_aw_bits_user = NastiRouter_io_slave_1_aw_bits_user;
  assign io_slaves_1_aw_bits_id = NastiRouter_io_slave_1_aw_bits_id;
  assign io_slaves_1_aw_bits_region = NastiRouter_io_slave_1_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = NastiRouter_io_slave_1_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = NastiRouter_io_slave_1_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = NastiRouter_io_slave_1_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = NastiRouter_io_slave_1_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = NastiRouter_io_slave_1_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = NastiRouter_io_slave_1_aw_bits_size;
  assign io_slaves_1_aw_bits_len = NastiRouter_io_slave_1_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = NastiRouter_io_slave_1_aw_bits_addr;
  assign io_slaves_1_aw_valid = NastiRouter_io_slave_1_aw_valid;
  assign io_masters_0_r_bits_user = NastiRouter_io_master_r_bits_user;
  assign io_masters_0_r_bits_id = NastiRouter_io_master_r_bits_id;
  assign io_masters_0_r_bits_last = NastiRouter_io_master_r_bits_last;
  assign io_masters_0_r_bits_data = NastiRouter_io_master_r_bits_data;
  assign io_masters_0_r_bits_resp = NastiRouter_io_master_r_bits_resp;
  assign io_masters_0_r_valid = NastiRouter_io_master_r_valid;
  assign io_masters_0_ar_ready = NastiRouter_io_master_ar_ready;
  assign io_masters_0_b_bits_user = NastiRouter_io_master_b_bits_user;
  assign io_masters_0_b_bits_id = NastiRouter_io_master_b_bits_id;
  assign io_masters_0_b_bits_resp = NastiRouter_io_master_b_bits_resp;
  assign io_masters_0_b_valid = NastiRouter_io_master_b_valid;
  assign io_masters_0_w_ready = NastiRouter_io_master_w_ready;
  assign io_masters_0_aw_ready = NastiRouter_io_master_aw_ready;
  NastiRouter_1 NastiRouter(.clk(clk), .reset(reset),
       .io_master_aw_ready( NastiRouter_io_master_aw_ready ),
       .io_master_aw_valid( io_masters_0_aw_valid ),
       .io_master_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_master_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_master_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_master_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_master_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_master_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_master_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_master_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_master_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_master_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_master_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_master_w_ready( NastiRouter_io_master_w_ready ),
       .io_master_w_valid( io_masters_0_w_valid ),
       .io_master_w_bits_data( io_masters_0_w_bits_data ),
       .io_master_w_bits_last( io_masters_0_w_bits_last ),
       .io_master_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_master_w_bits_user( io_masters_0_w_bits_user ),
       .io_master_b_ready( io_masters_0_b_ready ),
       .io_master_b_valid( NastiRouter_io_master_b_valid ),
       .io_master_b_bits_resp( NastiRouter_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiRouter_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiRouter_io_master_b_bits_user ),
       .io_master_ar_ready( NastiRouter_io_master_ar_ready ),
       .io_master_ar_valid( io_masters_0_ar_valid ),
       .io_master_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_master_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_master_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_master_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_master_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_master_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_master_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_master_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_master_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_master_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_master_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_master_r_ready( io_masters_0_r_ready ),
       .io_master_r_valid( NastiRouter_io_master_r_valid ),
       .io_master_r_bits_resp( NastiRouter_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiRouter_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiRouter_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiRouter_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiRouter_io_master_r_bits_user ),
       .io_slave_1_aw_ready( io_slaves_1_aw_ready ),
       .io_slave_1_aw_valid( NastiRouter_io_slave_1_aw_valid ),
       .io_slave_1_aw_bits_addr( NastiRouter_io_slave_1_aw_bits_addr ),
       .io_slave_1_aw_bits_len( NastiRouter_io_slave_1_aw_bits_len ),
       .io_slave_1_aw_bits_size( NastiRouter_io_slave_1_aw_bits_size ),
       .io_slave_1_aw_bits_burst( NastiRouter_io_slave_1_aw_bits_burst ),
       .io_slave_1_aw_bits_lock( NastiRouter_io_slave_1_aw_bits_lock ),
       .io_slave_1_aw_bits_cache( NastiRouter_io_slave_1_aw_bits_cache ),
       .io_slave_1_aw_bits_prot( NastiRouter_io_slave_1_aw_bits_prot ),
       .io_slave_1_aw_bits_qos( NastiRouter_io_slave_1_aw_bits_qos ),
       .io_slave_1_aw_bits_region( NastiRouter_io_slave_1_aw_bits_region ),
       .io_slave_1_aw_bits_id( NastiRouter_io_slave_1_aw_bits_id ),
       .io_slave_1_aw_bits_user( NastiRouter_io_slave_1_aw_bits_user ),
       .io_slave_1_w_ready( io_slaves_1_w_ready ),
       .io_slave_1_w_valid( NastiRouter_io_slave_1_w_valid ),
       .io_slave_1_w_bits_data( NastiRouter_io_slave_1_w_bits_data ),
       .io_slave_1_w_bits_last( NastiRouter_io_slave_1_w_bits_last ),
       .io_slave_1_w_bits_strb( NastiRouter_io_slave_1_w_bits_strb ),
       .io_slave_1_w_bits_user( NastiRouter_io_slave_1_w_bits_user ),
       .io_slave_1_b_ready( NastiRouter_io_slave_1_b_ready ),
       .io_slave_1_b_valid( io_slaves_1_b_valid ),
       .io_slave_1_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slave_1_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slave_1_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slave_1_ar_ready( io_slaves_1_ar_ready ),
       .io_slave_1_ar_valid( NastiRouter_io_slave_1_ar_valid ),
       .io_slave_1_ar_bits_addr( NastiRouter_io_slave_1_ar_bits_addr ),
       .io_slave_1_ar_bits_len( NastiRouter_io_slave_1_ar_bits_len ),
       .io_slave_1_ar_bits_size( NastiRouter_io_slave_1_ar_bits_size ),
       .io_slave_1_ar_bits_burst( NastiRouter_io_slave_1_ar_bits_burst ),
       .io_slave_1_ar_bits_lock( NastiRouter_io_slave_1_ar_bits_lock ),
       .io_slave_1_ar_bits_cache( NastiRouter_io_slave_1_ar_bits_cache ),
       .io_slave_1_ar_bits_prot( NastiRouter_io_slave_1_ar_bits_prot ),
       .io_slave_1_ar_bits_qos( NastiRouter_io_slave_1_ar_bits_qos ),
       .io_slave_1_ar_bits_region( NastiRouter_io_slave_1_ar_bits_region ),
       .io_slave_1_ar_bits_id( NastiRouter_io_slave_1_ar_bits_id ),
       .io_slave_1_ar_bits_user( NastiRouter_io_slave_1_ar_bits_user ),
       .io_slave_1_r_ready( NastiRouter_io_slave_1_r_ready ),
       .io_slave_1_r_valid( io_slaves_1_r_valid ),
       .io_slave_1_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slave_1_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slave_1_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slave_1_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slave_1_r_bits_user( io_slaves_1_r_bits_user ),
       .io_slave_0_aw_ready( io_slaves_0_aw_ready ),
       .io_slave_0_aw_valid( NastiRouter_io_slave_0_aw_valid ),
       .io_slave_0_aw_bits_addr( NastiRouter_io_slave_0_aw_bits_addr ),
       .io_slave_0_aw_bits_len( NastiRouter_io_slave_0_aw_bits_len ),
       .io_slave_0_aw_bits_size( NastiRouter_io_slave_0_aw_bits_size ),
       .io_slave_0_aw_bits_burst( NastiRouter_io_slave_0_aw_bits_burst ),
       .io_slave_0_aw_bits_lock( NastiRouter_io_slave_0_aw_bits_lock ),
       .io_slave_0_aw_bits_cache( NastiRouter_io_slave_0_aw_bits_cache ),
       .io_slave_0_aw_bits_prot( NastiRouter_io_slave_0_aw_bits_prot ),
       .io_slave_0_aw_bits_qos( NastiRouter_io_slave_0_aw_bits_qos ),
       .io_slave_0_aw_bits_region( NastiRouter_io_slave_0_aw_bits_region ),
       .io_slave_0_aw_bits_id( NastiRouter_io_slave_0_aw_bits_id ),
       .io_slave_0_aw_bits_user( NastiRouter_io_slave_0_aw_bits_user ),
       .io_slave_0_w_ready( io_slaves_0_w_ready ),
       .io_slave_0_w_valid( NastiRouter_io_slave_0_w_valid ),
       .io_slave_0_w_bits_data( NastiRouter_io_slave_0_w_bits_data ),
       .io_slave_0_w_bits_last( NastiRouter_io_slave_0_w_bits_last ),
       .io_slave_0_w_bits_strb( NastiRouter_io_slave_0_w_bits_strb ),
       .io_slave_0_w_bits_user( NastiRouter_io_slave_0_w_bits_user ),
       .io_slave_0_b_ready( NastiRouter_io_slave_0_b_ready ),
       .io_slave_0_b_valid( io_slaves_0_b_valid ),
       .io_slave_0_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slave_0_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slave_0_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slave_0_ar_ready( io_slaves_0_ar_ready ),
       .io_slave_0_ar_valid( NastiRouter_io_slave_0_ar_valid ),
       .io_slave_0_ar_bits_addr( NastiRouter_io_slave_0_ar_bits_addr ),
       .io_slave_0_ar_bits_len( NastiRouter_io_slave_0_ar_bits_len ),
       .io_slave_0_ar_bits_size( NastiRouter_io_slave_0_ar_bits_size ),
       .io_slave_0_ar_bits_burst( NastiRouter_io_slave_0_ar_bits_burst ),
       .io_slave_0_ar_bits_lock( NastiRouter_io_slave_0_ar_bits_lock ),
       .io_slave_0_ar_bits_cache( NastiRouter_io_slave_0_ar_bits_cache ),
       .io_slave_0_ar_bits_prot( NastiRouter_io_slave_0_ar_bits_prot ),
       .io_slave_0_ar_bits_qos( NastiRouter_io_slave_0_ar_bits_qos ),
       .io_slave_0_ar_bits_region( NastiRouter_io_slave_0_ar_bits_region ),
       .io_slave_0_ar_bits_id( NastiRouter_io_slave_0_ar_bits_id ),
       .io_slave_0_ar_bits_user( NastiRouter_io_slave_0_ar_bits_user ),
       .io_slave_0_r_ready( NastiRouter_io_slave_0_r_ready ),
       .io_slave_0_r_valid( io_slaves_0_r_valid ),
       .io_slave_0_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slave_0_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slave_0_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slave_0_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slave_0_r_bits_user( io_slaves_0_r_bits_user )
  );
endmodule

module NastiRecursiveInterconnect(input clk, input reset,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [4:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[4:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [4:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[4:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[4:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [4:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[4:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [4:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[4:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [4:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[4:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [4:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire xbar_io_masters_0_aw_ready;
  wire xbar_io_masters_0_w_ready;
  wire xbar_io_masters_0_b_valid;
  wire[1:0] xbar_io_masters_0_b_bits_resp;
  wire[4:0] xbar_io_masters_0_b_bits_id;
  wire xbar_io_masters_0_b_bits_user;
  wire xbar_io_masters_0_ar_ready;
  wire xbar_io_masters_0_r_valid;
  wire[1:0] xbar_io_masters_0_r_bits_resp;
  wire[63:0] xbar_io_masters_0_r_bits_data;
  wire xbar_io_masters_0_r_bits_last;
  wire[4:0] xbar_io_masters_0_r_bits_id;
  wire xbar_io_masters_0_r_bits_user;
  wire xbar_io_slaves_1_aw_valid;
  wire[31:0] xbar_io_slaves_1_aw_bits_addr;
  wire[7:0] xbar_io_slaves_1_aw_bits_len;
  wire[2:0] xbar_io_slaves_1_aw_bits_size;
  wire[1:0] xbar_io_slaves_1_aw_bits_burst;
  wire xbar_io_slaves_1_aw_bits_lock;
  wire[3:0] xbar_io_slaves_1_aw_bits_cache;
  wire[2:0] xbar_io_slaves_1_aw_bits_prot;
  wire[3:0] xbar_io_slaves_1_aw_bits_qos;
  wire[3:0] xbar_io_slaves_1_aw_bits_region;
  wire[4:0] xbar_io_slaves_1_aw_bits_id;
  wire xbar_io_slaves_1_aw_bits_user;
  wire xbar_io_slaves_1_w_valid;
  wire[63:0] xbar_io_slaves_1_w_bits_data;
  wire xbar_io_slaves_1_w_bits_last;
  wire[7:0] xbar_io_slaves_1_w_bits_strb;
  wire xbar_io_slaves_1_w_bits_user;
  wire xbar_io_slaves_1_b_ready;
  wire xbar_io_slaves_1_ar_valid;
  wire[31:0] xbar_io_slaves_1_ar_bits_addr;
  wire[7:0] xbar_io_slaves_1_ar_bits_len;
  wire[2:0] xbar_io_slaves_1_ar_bits_size;
  wire[1:0] xbar_io_slaves_1_ar_bits_burst;
  wire xbar_io_slaves_1_ar_bits_lock;
  wire[3:0] xbar_io_slaves_1_ar_bits_cache;
  wire[2:0] xbar_io_slaves_1_ar_bits_prot;
  wire[3:0] xbar_io_slaves_1_ar_bits_qos;
  wire[3:0] xbar_io_slaves_1_ar_bits_region;
  wire[4:0] xbar_io_slaves_1_ar_bits_id;
  wire xbar_io_slaves_1_ar_bits_user;
  wire xbar_io_slaves_1_r_ready;
  wire xbar_io_slaves_0_aw_valid;
  wire[31:0] xbar_io_slaves_0_aw_bits_addr;
  wire[7:0] xbar_io_slaves_0_aw_bits_len;
  wire[2:0] xbar_io_slaves_0_aw_bits_size;
  wire[1:0] xbar_io_slaves_0_aw_bits_burst;
  wire xbar_io_slaves_0_aw_bits_lock;
  wire[3:0] xbar_io_slaves_0_aw_bits_cache;
  wire[2:0] xbar_io_slaves_0_aw_bits_prot;
  wire[3:0] xbar_io_slaves_0_aw_bits_qos;
  wire[3:0] xbar_io_slaves_0_aw_bits_region;
  wire[4:0] xbar_io_slaves_0_aw_bits_id;
  wire xbar_io_slaves_0_aw_bits_user;
  wire xbar_io_slaves_0_w_valid;
  wire[63:0] xbar_io_slaves_0_w_bits_data;
  wire xbar_io_slaves_0_w_bits_last;
  wire[7:0] xbar_io_slaves_0_w_bits_strb;
  wire xbar_io_slaves_0_w_bits_user;
  wire xbar_io_slaves_0_b_ready;
  wire xbar_io_slaves_0_ar_valid;
  wire[31:0] xbar_io_slaves_0_ar_bits_addr;
  wire[7:0] xbar_io_slaves_0_ar_bits_len;
  wire[2:0] xbar_io_slaves_0_ar_bits_size;
  wire[1:0] xbar_io_slaves_0_ar_bits_burst;
  wire xbar_io_slaves_0_ar_bits_lock;
  wire[3:0] xbar_io_slaves_0_ar_bits_cache;
  wire[2:0] xbar_io_slaves_0_ar_bits_prot;
  wire[3:0] xbar_io_slaves_0_ar_bits_qos;
  wire[3:0] xbar_io_slaves_0_ar_bits_region;
  wire[4:0] xbar_io_slaves_0_ar_bits_id;
  wire xbar_io_slaves_0_ar_bits_user;
  wire xbar_io_slaves_0_r_ready;


  assign io_slaves_0_r_ready = xbar_io_slaves_0_r_ready;
  assign io_slaves_0_ar_bits_user = xbar_io_slaves_0_ar_bits_user;
  assign io_slaves_0_ar_bits_id = xbar_io_slaves_0_ar_bits_id;
  assign io_slaves_0_ar_bits_region = xbar_io_slaves_0_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = xbar_io_slaves_0_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = xbar_io_slaves_0_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = xbar_io_slaves_0_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = xbar_io_slaves_0_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = xbar_io_slaves_0_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = xbar_io_slaves_0_ar_bits_size;
  assign io_slaves_0_ar_bits_len = xbar_io_slaves_0_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = xbar_io_slaves_0_ar_bits_addr;
  assign io_slaves_0_ar_valid = xbar_io_slaves_0_ar_valid;
  assign io_slaves_0_b_ready = xbar_io_slaves_0_b_ready;
  assign io_slaves_0_w_bits_user = xbar_io_slaves_0_w_bits_user;
  assign io_slaves_0_w_bits_strb = xbar_io_slaves_0_w_bits_strb;
  assign io_slaves_0_w_bits_last = xbar_io_slaves_0_w_bits_last;
  assign io_slaves_0_w_bits_data = xbar_io_slaves_0_w_bits_data;
  assign io_slaves_0_w_valid = xbar_io_slaves_0_w_valid;
  assign io_slaves_0_aw_bits_user = xbar_io_slaves_0_aw_bits_user;
  assign io_slaves_0_aw_bits_id = xbar_io_slaves_0_aw_bits_id;
  assign io_slaves_0_aw_bits_region = xbar_io_slaves_0_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = xbar_io_slaves_0_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = xbar_io_slaves_0_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = xbar_io_slaves_0_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = xbar_io_slaves_0_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = xbar_io_slaves_0_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = xbar_io_slaves_0_aw_bits_size;
  assign io_slaves_0_aw_bits_len = xbar_io_slaves_0_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = xbar_io_slaves_0_aw_bits_addr;
  assign io_slaves_0_aw_valid = xbar_io_slaves_0_aw_valid;
  assign io_slaves_1_r_ready = xbar_io_slaves_1_r_ready;
  assign io_slaves_1_ar_bits_user = xbar_io_slaves_1_ar_bits_user;
  assign io_slaves_1_ar_bits_id = xbar_io_slaves_1_ar_bits_id;
  assign io_slaves_1_ar_bits_region = xbar_io_slaves_1_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = xbar_io_slaves_1_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = xbar_io_slaves_1_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = xbar_io_slaves_1_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = xbar_io_slaves_1_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = xbar_io_slaves_1_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = xbar_io_slaves_1_ar_bits_size;
  assign io_slaves_1_ar_bits_len = xbar_io_slaves_1_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = xbar_io_slaves_1_ar_bits_addr;
  assign io_slaves_1_ar_valid = xbar_io_slaves_1_ar_valid;
  assign io_slaves_1_b_ready = xbar_io_slaves_1_b_ready;
  assign io_slaves_1_w_bits_user = xbar_io_slaves_1_w_bits_user;
  assign io_slaves_1_w_bits_strb = xbar_io_slaves_1_w_bits_strb;
  assign io_slaves_1_w_bits_last = xbar_io_slaves_1_w_bits_last;
  assign io_slaves_1_w_bits_data = xbar_io_slaves_1_w_bits_data;
  assign io_slaves_1_w_valid = xbar_io_slaves_1_w_valid;
  assign io_slaves_1_aw_bits_user = xbar_io_slaves_1_aw_bits_user;
  assign io_slaves_1_aw_bits_id = xbar_io_slaves_1_aw_bits_id;
  assign io_slaves_1_aw_bits_region = xbar_io_slaves_1_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = xbar_io_slaves_1_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = xbar_io_slaves_1_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = xbar_io_slaves_1_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = xbar_io_slaves_1_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = xbar_io_slaves_1_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = xbar_io_slaves_1_aw_bits_size;
  assign io_slaves_1_aw_bits_len = xbar_io_slaves_1_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = xbar_io_slaves_1_aw_bits_addr;
  assign io_slaves_1_aw_valid = xbar_io_slaves_1_aw_valid;
  assign io_masters_0_r_bits_user = xbar_io_masters_0_r_bits_user;
  assign io_masters_0_r_bits_id = xbar_io_masters_0_r_bits_id;
  assign io_masters_0_r_bits_last = xbar_io_masters_0_r_bits_last;
  assign io_masters_0_r_bits_data = xbar_io_masters_0_r_bits_data;
  assign io_masters_0_r_bits_resp = xbar_io_masters_0_r_bits_resp;
  assign io_masters_0_r_valid = xbar_io_masters_0_r_valid;
  assign io_masters_0_ar_ready = xbar_io_masters_0_ar_ready;
  assign io_masters_0_b_bits_user = xbar_io_masters_0_b_bits_user;
  assign io_masters_0_b_bits_id = xbar_io_masters_0_b_bits_id;
  assign io_masters_0_b_bits_resp = xbar_io_masters_0_b_bits_resp;
  assign io_masters_0_b_valid = xbar_io_masters_0_b_valid;
  assign io_masters_0_w_ready = xbar_io_masters_0_w_ready;
  assign io_masters_0_aw_ready = xbar_io_masters_0_aw_ready;
  NastiCrossbar_1 xbar(.clk(clk), .reset(reset),
       .io_masters_0_aw_ready( xbar_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( io_masters_0_aw_valid ),
       .io_masters_0_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_masters_0_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_masters_0_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_masters_0_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_masters_0_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_masters_0_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_masters_0_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_masters_0_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_masters_0_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_masters_0_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_masters_0_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_masters_0_w_ready( xbar_io_masters_0_w_ready ),
       .io_masters_0_w_valid( io_masters_0_w_valid ),
       .io_masters_0_w_bits_data( io_masters_0_w_bits_data ),
       .io_masters_0_w_bits_last( io_masters_0_w_bits_last ),
       .io_masters_0_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_masters_0_w_bits_user( io_masters_0_w_bits_user ),
       .io_masters_0_b_ready( io_masters_0_b_ready ),
       .io_masters_0_b_valid( xbar_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( xbar_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( xbar_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( xbar_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( xbar_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( io_masters_0_ar_valid ),
       .io_masters_0_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_masters_0_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_masters_0_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_masters_0_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_masters_0_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_masters_0_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_masters_0_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_masters_0_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_masters_0_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_masters_0_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_masters_0_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_masters_0_r_ready( io_masters_0_r_ready ),
       .io_masters_0_r_valid( xbar_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( xbar_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( xbar_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( xbar_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( xbar_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( xbar_io_masters_0_r_bits_user ),
       .io_slaves_1_aw_ready( io_slaves_1_aw_ready ),
       .io_slaves_1_aw_valid( xbar_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( xbar_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( xbar_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( xbar_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( xbar_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( xbar_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( xbar_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( xbar_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( xbar_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( xbar_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( xbar_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( xbar_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( io_slaves_1_w_ready ),
       .io_slaves_1_w_valid( xbar_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( xbar_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( xbar_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( xbar_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( xbar_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( xbar_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( io_slaves_1_b_valid ),
       .io_slaves_1_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slaves_1_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slaves_1_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slaves_1_ar_ready( io_slaves_1_ar_ready ),
       .io_slaves_1_ar_valid( xbar_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( xbar_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( xbar_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( xbar_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( xbar_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( xbar_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( xbar_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( xbar_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( xbar_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( xbar_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( xbar_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( xbar_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( xbar_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( io_slaves_1_r_valid ),
       .io_slaves_1_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slaves_1_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slaves_1_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slaves_1_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slaves_1_r_bits_user( io_slaves_1_r_bits_user ),
       .io_slaves_0_aw_ready( io_slaves_0_aw_ready ),
       .io_slaves_0_aw_valid( xbar_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( xbar_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( xbar_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( xbar_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( xbar_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( xbar_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( xbar_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( xbar_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( xbar_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( xbar_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( xbar_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( xbar_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_slaves_0_w_ready ),
       .io_slaves_0_w_valid( xbar_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( xbar_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( xbar_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( xbar_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( xbar_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( xbar_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_slaves_0_b_valid ),
       .io_slaves_0_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slaves_0_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slaves_0_ar_ready( io_slaves_0_ar_ready ),
       .io_slaves_0_ar_valid( xbar_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( xbar_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( xbar_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( xbar_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( xbar_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( xbar_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( xbar_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( xbar_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( xbar_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( xbar_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( xbar_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( xbar_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( xbar_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_slaves_0_r_valid ),
       .io_slaves_0_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slaves_0_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slaves_0_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slaves_0_r_bits_user( io_slaves_0_r_bits_user )
  );
endmodule

module NastiRecursiveInterconnect_1(input clk, input reset,
    output io_masters_1_aw_ready,
    input  io_masters_1_aw_valid,
    input [31:0] io_masters_1_aw_bits_addr,
    input [7:0] io_masters_1_aw_bits_len,
    input [2:0] io_masters_1_aw_bits_size,
    input [1:0] io_masters_1_aw_bits_burst,
    input  io_masters_1_aw_bits_lock,
    input [3:0] io_masters_1_aw_bits_cache,
    input [2:0] io_masters_1_aw_bits_prot,
    input [3:0] io_masters_1_aw_bits_qos,
    input [3:0] io_masters_1_aw_bits_region,
    input [4:0] io_masters_1_aw_bits_id,
    input  io_masters_1_aw_bits_user,
    output io_masters_1_w_ready,
    input  io_masters_1_w_valid,
    input [63:0] io_masters_1_w_bits_data,
    input  io_masters_1_w_bits_last,
    input [7:0] io_masters_1_w_bits_strb,
    input  io_masters_1_w_bits_user,
    input  io_masters_1_b_ready,
    output io_masters_1_b_valid,
    output[1:0] io_masters_1_b_bits_resp,
    output[4:0] io_masters_1_b_bits_id,
    output io_masters_1_b_bits_user,
    output io_masters_1_ar_ready,
    input  io_masters_1_ar_valid,
    input [31:0] io_masters_1_ar_bits_addr,
    input [7:0] io_masters_1_ar_bits_len,
    input [2:0] io_masters_1_ar_bits_size,
    input [1:0] io_masters_1_ar_bits_burst,
    input  io_masters_1_ar_bits_lock,
    input [3:0] io_masters_1_ar_bits_cache,
    input [2:0] io_masters_1_ar_bits_prot,
    input [3:0] io_masters_1_ar_bits_qos,
    input [3:0] io_masters_1_ar_bits_region,
    input [4:0] io_masters_1_ar_bits_id,
    input  io_masters_1_ar_bits_user,
    input  io_masters_1_r_ready,
    output io_masters_1_r_valid,
    output[1:0] io_masters_1_r_bits_resp,
    output[63:0] io_masters_1_r_bits_data,
    output io_masters_1_r_bits_last,
    output[4:0] io_masters_1_r_bits_id,
    output io_masters_1_r_bits_user,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [4:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[4:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [4:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[4:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_3_aw_ready,
    output io_slaves_3_aw_valid,
    output[31:0] io_slaves_3_aw_bits_addr,
    output[7:0] io_slaves_3_aw_bits_len,
    output[2:0] io_slaves_3_aw_bits_size,
    output[1:0] io_slaves_3_aw_bits_burst,
    output io_slaves_3_aw_bits_lock,
    output[3:0] io_slaves_3_aw_bits_cache,
    output[2:0] io_slaves_3_aw_bits_prot,
    output[3:0] io_slaves_3_aw_bits_qos,
    output[3:0] io_slaves_3_aw_bits_region,
    output[4:0] io_slaves_3_aw_bits_id,
    output io_slaves_3_aw_bits_user,
    input  io_slaves_3_w_ready,
    output io_slaves_3_w_valid,
    output[63:0] io_slaves_3_w_bits_data,
    output io_slaves_3_w_bits_last,
    output[7:0] io_slaves_3_w_bits_strb,
    output io_slaves_3_w_bits_user,
    output io_slaves_3_b_ready,
    input  io_slaves_3_b_valid,
    input [1:0] io_slaves_3_b_bits_resp,
    input [4:0] io_slaves_3_b_bits_id,
    input  io_slaves_3_b_bits_user,
    input  io_slaves_3_ar_ready,
    output io_slaves_3_ar_valid,
    output[31:0] io_slaves_3_ar_bits_addr,
    output[7:0] io_slaves_3_ar_bits_len,
    output[2:0] io_slaves_3_ar_bits_size,
    output[1:0] io_slaves_3_ar_bits_burst,
    output io_slaves_3_ar_bits_lock,
    output[3:0] io_slaves_3_ar_bits_cache,
    output[2:0] io_slaves_3_ar_bits_prot,
    output[3:0] io_slaves_3_ar_bits_qos,
    output[3:0] io_slaves_3_ar_bits_region,
    output[4:0] io_slaves_3_ar_bits_id,
    output io_slaves_3_ar_bits_user,
    output io_slaves_3_r_ready,
    input  io_slaves_3_r_valid,
    input [1:0] io_slaves_3_r_bits_resp,
    input [63:0] io_slaves_3_r_bits_data,
    input  io_slaves_3_r_bits_last,
    input [4:0] io_slaves_3_r_bits_id,
    input  io_slaves_3_r_bits_user,
    input  io_slaves_2_aw_ready,
    output io_slaves_2_aw_valid,
    output[31:0] io_slaves_2_aw_bits_addr,
    output[7:0] io_slaves_2_aw_bits_len,
    output[2:0] io_slaves_2_aw_bits_size,
    output[1:0] io_slaves_2_aw_bits_burst,
    output io_slaves_2_aw_bits_lock,
    output[3:0] io_slaves_2_aw_bits_cache,
    output[2:0] io_slaves_2_aw_bits_prot,
    output[3:0] io_slaves_2_aw_bits_qos,
    output[3:0] io_slaves_2_aw_bits_region,
    output[4:0] io_slaves_2_aw_bits_id,
    output io_slaves_2_aw_bits_user,
    input  io_slaves_2_w_ready,
    output io_slaves_2_w_valid,
    output[63:0] io_slaves_2_w_bits_data,
    output io_slaves_2_w_bits_last,
    output[7:0] io_slaves_2_w_bits_strb,
    output io_slaves_2_w_bits_user,
    output io_slaves_2_b_ready,
    input  io_slaves_2_b_valid,
    input [1:0] io_slaves_2_b_bits_resp,
    input [4:0] io_slaves_2_b_bits_id,
    input  io_slaves_2_b_bits_user,
    input  io_slaves_2_ar_ready,
    output io_slaves_2_ar_valid,
    output[31:0] io_slaves_2_ar_bits_addr,
    output[7:0] io_slaves_2_ar_bits_len,
    output[2:0] io_slaves_2_ar_bits_size,
    output[1:0] io_slaves_2_ar_bits_burst,
    output io_slaves_2_ar_bits_lock,
    output[3:0] io_slaves_2_ar_bits_cache,
    output[2:0] io_slaves_2_ar_bits_prot,
    output[3:0] io_slaves_2_ar_bits_qos,
    output[3:0] io_slaves_2_ar_bits_region,
    output[4:0] io_slaves_2_ar_bits_id,
    output io_slaves_2_ar_bits_user,
    output io_slaves_2_r_ready,
    input  io_slaves_2_r_valid,
    input [1:0] io_slaves_2_r_bits_resp,
    input [63:0] io_slaves_2_r_bits_data,
    input  io_slaves_2_r_bits_last,
    input [4:0] io_slaves_2_r_bits_id,
    input  io_slaves_2_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[4:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [4:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[4:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [4:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[4:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [4:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[4:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [4:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire NastiMultiChannelRouter_io_master_aw_ready;
  wire NastiMultiChannelRouter_io_master_w_ready;
  wire NastiMultiChannelRouter_io_master_b_valid;
  wire[1:0] NastiMultiChannelRouter_io_master_b_bits_resp;
  wire[4:0] NastiMultiChannelRouter_io_master_b_bits_id;
  wire NastiMultiChannelRouter_io_master_b_bits_user;
  wire NastiMultiChannelRouter_io_master_ar_ready;
  wire NastiMultiChannelRouter_io_master_r_valid;
  wire[1:0] NastiMultiChannelRouter_io_master_r_bits_resp;
  wire[63:0] NastiMultiChannelRouter_io_master_r_bits_data;
  wire NastiMultiChannelRouter_io_master_r_bits_last;
  wire[4:0] NastiMultiChannelRouter_io_master_r_bits_id;
  wire NastiMultiChannelRouter_io_master_r_bits_user;
  wire NastiMultiChannelRouter_io_slaves_0_aw_valid;
  wire[31:0] NastiMultiChannelRouter_io_slaves_0_aw_bits_addr;
  wire[7:0] NastiMultiChannelRouter_io_slaves_0_aw_bits_len;
  wire[2:0] NastiMultiChannelRouter_io_slaves_0_aw_bits_size;
  wire[1:0] NastiMultiChannelRouter_io_slaves_0_aw_bits_burst;
  wire NastiMultiChannelRouter_io_slaves_0_aw_bits_lock;
  wire[3:0] NastiMultiChannelRouter_io_slaves_0_aw_bits_cache;
  wire[2:0] NastiMultiChannelRouter_io_slaves_0_aw_bits_prot;
  wire[3:0] NastiMultiChannelRouter_io_slaves_0_aw_bits_qos;
  wire[3:0] NastiMultiChannelRouter_io_slaves_0_aw_bits_region;
  wire[4:0] NastiMultiChannelRouter_io_slaves_0_aw_bits_id;
  wire NastiMultiChannelRouter_io_slaves_0_aw_bits_user;
  wire NastiMultiChannelRouter_io_slaves_0_w_valid;
  wire[63:0] NastiMultiChannelRouter_io_slaves_0_w_bits_data;
  wire NastiMultiChannelRouter_io_slaves_0_w_bits_last;
  wire[7:0] NastiMultiChannelRouter_io_slaves_0_w_bits_strb;
  wire NastiMultiChannelRouter_io_slaves_0_w_bits_user;
  wire NastiMultiChannelRouter_io_slaves_0_b_ready;
  wire NastiMultiChannelRouter_io_slaves_0_ar_valid;
  wire[31:0] NastiMultiChannelRouter_io_slaves_0_ar_bits_addr;
  wire[7:0] NastiMultiChannelRouter_io_slaves_0_ar_bits_len;
  wire[2:0] NastiMultiChannelRouter_io_slaves_0_ar_bits_size;
  wire[1:0] NastiMultiChannelRouter_io_slaves_0_ar_bits_burst;
  wire NastiMultiChannelRouter_io_slaves_0_ar_bits_lock;
  wire[3:0] NastiMultiChannelRouter_io_slaves_0_ar_bits_cache;
  wire[2:0] NastiMultiChannelRouter_io_slaves_0_ar_bits_prot;
  wire[3:0] NastiMultiChannelRouter_io_slaves_0_ar_bits_qos;
  wire[3:0] NastiMultiChannelRouter_io_slaves_0_ar_bits_region;
  wire[4:0] NastiMultiChannelRouter_io_slaves_0_ar_bits_id;
  wire NastiMultiChannelRouter_io_slaves_0_ar_bits_user;
  wire NastiMultiChannelRouter_io_slaves_0_r_ready;
  wire xbar_io_masters_1_aw_ready;
  wire xbar_io_masters_1_w_ready;
  wire xbar_io_masters_1_b_valid;
  wire[1:0] xbar_io_masters_1_b_bits_resp;
  wire[4:0] xbar_io_masters_1_b_bits_id;
  wire xbar_io_masters_1_b_bits_user;
  wire xbar_io_masters_1_ar_ready;
  wire xbar_io_masters_1_r_valid;
  wire[1:0] xbar_io_masters_1_r_bits_resp;
  wire[63:0] xbar_io_masters_1_r_bits_data;
  wire xbar_io_masters_1_r_bits_last;
  wire[4:0] xbar_io_masters_1_r_bits_id;
  wire xbar_io_masters_1_r_bits_user;
  wire xbar_io_masters_0_aw_ready;
  wire xbar_io_masters_0_w_ready;
  wire xbar_io_masters_0_b_valid;
  wire[1:0] xbar_io_masters_0_b_bits_resp;
  wire[4:0] xbar_io_masters_0_b_bits_id;
  wire xbar_io_masters_0_b_bits_user;
  wire xbar_io_masters_0_ar_ready;
  wire xbar_io_masters_0_r_valid;
  wire[1:0] xbar_io_masters_0_r_bits_resp;
  wire[63:0] xbar_io_masters_0_r_bits_data;
  wire xbar_io_masters_0_r_bits_last;
  wire[4:0] xbar_io_masters_0_r_bits_id;
  wire xbar_io_masters_0_r_bits_user;
  wire xbar_io_slaves_2_aw_valid;
  wire[31:0] xbar_io_slaves_2_aw_bits_addr;
  wire[7:0] xbar_io_slaves_2_aw_bits_len;
  wire[2:0] xbar_io_slaves_2_aw_bits_size;
  wire[1:0] xbar_io_slaves_2_aw_bits_burst;
  wire xbar_io_slaves_2_aw_bits_lock;
  wire[3:0] xbar_io_slaves_2_aw_bits_cache;
  wire[2:0] xbar_io_slaves_2_aw_bits_prot;
  wire[3:0] xbar_io_slaves_2_aw_bits_qos;
  wire[3:0] xbar_io_slaves_2_aw_bits_region;
  wire[4:0] xbar_io_slaves_2_aw_bits_id;
  wire xbar_io_slaves_2_aw_bits_user;
  wire xbar_io_slaves_2_w_valid;
  wire[63:0] xbar_io_slaves_2_w_bits_data;
  wire xbar_io_slaves_2_w_bits_last;
  wire[7:0] xbar_io_slaves_2_w_bits_strb;
  wire xbar_io_slaves_2_w_bits_user;
  wire xbar_io_slaves_2_b_ready;
  wire xbar_io_slaves_2_ar_valid;
  wire[31:0] xbar_io_slaves_2_ar_bits_addr;
  wire[7:0] xbar_io_slaves_2_ar_bits_len;
  wire[2:0] xbar_io_slaves_2_ar_bits_size;
  wire[1:0] xbar_io_slaves_2_ar_bits_burst;
  wire xbar_io_slaves_2_ar_bits_lock;
  wire[3:0] xbar_io_slaves_2_ar_bits_cache;
  wire[2:0] xbar_io_slaves_2_ar_bits_prot;
  wire[3:0] xbar_io_slaves_2_ar_bits_qos;
  wire[3:0] xbar_io_slaves_2_ar_bits_region;
  wire[4:0] xbar_io_slaves_2_ar_bits_id;
  wire xbar_io_slaves_2_ar_bits_user;
  wire xbar_io_slaves_2_r_ready;
  wire xbar_io_slaves_1_aw_valid;
  wire[31:0] xbar_io_slaves_1_aw_bits_addr;
  wire[7:0] xbar_io_slaves_1_aw_bits_len;
  wire[2:0] xbar_io_slaves_1_aw_bits_size;
  wire[1:0] xbar_io_slaves_1_aw_bits_burst;
  wire xbar_io_slaves_1_aw_bits_lock;
  wire[3:0] xbar_io_slaves_1_aw_bits_cache;
  wire[2:0] xbar_io_slaves_1_aw_bits_prot;
  wire[3:0] xbar_io_slaves_1_aw_bits_qos;
  wire[3:0] xbar_io_slaves_1_aw_bits_region;
  wire[4:0] xbar_io_slaves_1_aw_bits_id;
  wire xbar_io_slaves_1_aw_bits_user;
  wire xbar_io_slaves_1_w_valid;
  wire[63:0] xbar_io_slaves_1_w_bits_data;
  wire xbar_io_slaves_1_w_bits_last;
  wire[7:0] xbar_io_slaves_1_w_bits_strb;
  wire xbar_io_slaves_1_w_bits_user;
  wire xbar_io_slaves_1_b_ready;
  wire xbar_io_slaves_1_ar_valid;
  wire[31:0] xbar_io_slaves_1_ar_bits_addr;
  wire[7:0] xbar_io_slaves_1_ar_bits_len;
  wire[2:0] xbar_io_slaves_1_ar_bits_size;
  wire[1:0] xbar_io_slaves_1_ar_bits_burst;
  wire xbar_io_slaves_1_ar_bits_lock;
  wire[3:0] xbar_io_slaves_1_ar_bits_cache;
  wire[2:0] xbar_io_slaves_1_ar_bits_prot;
  wire[3:0] xbar_io_slaves_1_ar_bits_qos;
  wire[3:0] xbar_io_slaves_1_ar_bits_region;
  wire[4:0] xbar_io_slaves_1_ar_bits_id;
  wire xbar_io_slaves_1_ar_bits_user;
  wire xbar_io_slaves_1_r_ready;
  wire xbar_io_slaves_0_aw_valid;
  wire[31:0] xbar_io_slaves_0_aw_bits_addr;
  wire[7:0] xbar_io_slaves_0_aw_bits_len;
  wire[2:0] xbar_io_slaves_0_aw_bits_size;
  wire[1:0] xbar_io_slaves_0_aw_bits_burst;
  wire xbar_io_slaves_0_aw_bits_lock;
  wire[3:0] xbar_io_slaves_0_aw_bits_cache;
  wire[2:0] xbar_io_slaves_0_aw_bits_prot;
  wire[3:0] xbar_io_slaves_0_aw_bits_qos;
  wire[3:0] xbar_io_slaves_0_aw_bits_region;
  wire[4:0] xbar_io_slaves_0_aw_bits_id;
  wire xbar_io_slaves_0_aw_bits_user;
  wire xbar_io_slaves_0_w_valid;
  wire[63:0] xbar_io_slaves_0_w_bits_data;
  wire xbar_io_slaves_0_w_bits_last;
  wire[7:0] xbar_io_slaves_0_w_bits_strb;
  wire xbar_io_slaves_0_w_bits_user;
  wire xbar_io_slaves_0_b_ready;
  wire xbar_io_slaves_0_ar_valid;
  wire[31:0] xbar_io_slaves_0_ar_bits_addr;
  wire[7:0] xbar_io_slaves_0_ar_bits_len;
  wire[2:0] xbar_io_slaves_0_ar_bits_size;
  wire[1:0] xbar_io_slaves_0_ar_bits_burst;
  wire xbar_io_slaves_0_ar_bits_lock;
  wire[3:0] xbar_io_slaves_0_ar_bits_cache;
  wire[2:0] xbar_io_slaves_0_ar_bits_prot;
  wire[3:0] xbar_io_slaves_0_ar_bits_qos;
  wire[3:0] xbar_io_slaves_0_ar_bits_region;
  wire[4:0] xbar_io_slaves_0_ar_bits_id;
  wire xbar_io_slaves_0_ar_bits_user;
  wire xbar_io_slaves_0_r_ready;
  wire NastiRecursiveInterconnect_io_masters_0_aw_ready;
  wire NastiRecursiveInterconnect_io_masters_0_w_ready;
  wire NastiRecursiveInterconnect_io_masters_0_b_valid;
  wire[1:0] NastiRecursiveInterconnect_io_masters_0_b_bits_resp;
  wire[4:0] NastiRecursiveInterconnect_io_masters_0_b_bits_id;
  wire NastiRecursiveInterconnect_io_masters_0_b_bits_user;
  wire NastiRecursiveInterconnect_io_masters_0_ar_ready;
  wire NastiRecursiveInterconnect_io_masters_0_r_valid;
  wire[1:0] NastiRecursiveInterconnect_io_masters_0_r_bits_resp;
  wire[63:0] NastiRecursiveInterconnect_io_masters_0_r_bits_data;
  wire NastiRecursiveInterconnect_io_masters_0_r_bits_last;
  wire[4:0] NastiRecursiveInterconnect_io_masters_0_r_bits_id;
  wire NastiRecursiveInterconnect_io_masters_0_r_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_aw_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_1_aw_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_region;
  wire[4:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_1_aw_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_w_valid;
  wire[63:0] NastiRecursiveInterconnect_io_slaves_1_w_bits_data;
  wire NastiRecursiveInterconnect_io_slaves_1_w_bits_last;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_1_w_bits_strb;
  wire NastiRecursiveInterconnect_io_slaves_1_w_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_b_ready;
  wire NastiRecursiveInterconnect_io_slaves_1_ar_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_1_ar_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_region;
  wire[4:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_1_ar_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_r_ready;
  wire NastiRecursiveInterconnect_io_slaves_0_aw_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_0_aw_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_region;
  wire[4:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_0_aw_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_0_w_valid;
  wire[63:0] NastiRecursiveInterconnect_io_slaves_0_w_bits_data;
  wire NastiRecursiveInterconnect_io_slaves_0_w_bits_last;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_0_w_bits_strb;
  wire NastiRecursiveInterconnect_io_slaves_0_w_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_0_b_ready;
  wire NastiRecursiveInterconnect_io_slaves_0_ar_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_0_ar_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_region;
  wire[4:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_0_ar_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_0_r_ready;


  assign io_slaves_0_r_ready = NastiMultiChannelRouter_io_slaves_0_r_ready;
  assign io_slaves_0_ar_bits_user = NastiMultiChannelRouter_io_slaves_0_ar_bits_user;
  assign io_slaves_0_ar_bits_id = NastiMultiChannelRouter_io_slaves_0_ar_bits_id;
  assign io_slaves_0_ar_bits_region = NastiMultiChannelRouter_io_slaves_0_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = NastiMultiChannelRouter_io_slaves_0_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = NastiMultiChannelRouter_io_slaves_0_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = NastiMultiChannelRouter_io_slaves_0_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = NastiMultiChannelRouter_io_slaves_0_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = NastiMultiChannelRouter_io_slaves_0_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = NastiMultiChannelRouter_io_slaves_0_ar_bits_size;
  assign io_slaves_0_ar_bits_len = NastiMultiChannelRouter_io_slaves_0_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = NastiMultiChannelRouter_io_slaves_0_ar_bits_addr;
  assign io_slaves_0_ar_valid = NastiMultiChannelRouter_io_slaves_0_ar_valid;
  assign io_slaves_0_b_ready = NastiMultiChannelRouter_io_slaves_0_b_ready;
  assign io_slaves_0_w_bits_user = NastiMultiChannelRouter_io_slaves_0_w_bits_user;
  assign io_slaves_0_w_bits_strb = NastiMultiChannelRouter_io_slaves_0_w_bits_strb;
  assign io_slaves_0_w_bits_last = NastiMultiChannelRouter_io_slaves_0_w_bits_last;
  assign io_slaves_0_w_bits_data = NastiMultiChannelRouter_io_slaves_0_w_bits_data;
  assign io_slaves_0_w_valid = NastiMultiChannelRouter_io_slaves_0_w_valid;
  assign io_slaves_0_aw_bits_user = NastiMultiChannelRouter_io_slaves_0_aw_bits_user;
  assign io_slaves_0_aw_bits_id = NastiMultiChannelRouter_io_slaves_0_aw_bits_id;
  assign io_slaves_0_aw_bits_region = NastiMultiChannelRouter_io_slaves_0_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = NastiMultiChannelRouter_io_slaves_0_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = NastiMultiChannelRouter_io_slaves_0_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = NastiMultiChannelRouter_io_slaves_0_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = NastiMultiChannelRouter_io_slaves_0_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = NastiMultiChannelRouter_io_slaves_0_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = NastiMultiChannelRouter_io_slaves_0_aw_bits_size;
  assign io_slaves_0_aw_bits_len = NastiMultiChannelRouter_io_slaves_0_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = NastiMultiChannelRouter_io_slaves_0_aw_bits_addr;
  assign io_slaves_0_aw_valid = NastiMultiChannelRouter_io_slaves_0_aw_valid;
  assign io_slaves_1_r_ready = NastiRecursiveInterconnect_io_slaves_0_r_ready;
  assign io_slaves_1_ar_bits_user = NastiRecursiveInterconnect_io_slaves_0_ar_bits_user;
  assign io_slaves_1_ar_bits_id = NastiRecursiveInterconnect_io_slaves_0_ar_bits_id;
  assign io_slaves_1_ar_bits_region = NastiRecursiveInterconnect_io_slaves_0_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = NastiRecursiveInterconnect_io_slaves_0_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = NastiRecursiveInterconnect_io_slaves_0_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = NastiRecursiveInterconnect_io_slaves_0_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = NastiRecursiveInterconnect_io_slaves_0_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = NastiRecursiveInterconnect_io_slaves_0_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = NastiRecursiveInterconnect_io_slaves_0_ar_bits_size;
  assign io_slaves_1_ar_bits_len = NastiRecursiveInterconnect_io_slaves_0_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = NastiRecursiveInterconnect_io_slaves_0_ar_bits_addr;
  assign io_slaves_1_ar_valid = NastiRecursiveInterconnect_io_slaves_0_ar_valid;
  assign io_slaves_1_b_ready = NastiRecursiveInterconnect_io_slaves_0_b_ready;
  assign io_slaves_1_w_bits_user = NastiRecursiveInterconnect_io_slaves_0_w_bits_user;
  assign io_slaves_1_w_bits_strb = NastiRecursiveInterconnect_io_slaves_0_w_bits_strb;
  assign io_slaves_1_w_bits_last = NastiRecursiveInterconnect_io_slaves_0_w_bits_last;
  assign io_slaves_1_w_bits_data = NastiRecursiveInterconnect_io_slaves_0_w_bits_data;
  assign io_slaves_1_w_valid = NastiRecursiveInterconnect_io_slaves_0_w_valid;
  assign io_slaves_1_aw_bits_user = NastiRecursiveInterconnect_io_slaves_0_aw_bits_user;
  assign io_slaves_1_aw_bits_id = NastiRecursiveInterconnect_io_slaves_0_aw_bits_id;
  assign io_slaves_1_aw_bits_region = NastiRecursiveInterconnect_io_slaves_0_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = NastiRecursiveInterconnect_io_slaves_0_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = NastiRecursiveInterconnect_io_slaves_0_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = NastiRecursiveInterconnect_io_slaves_0_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = NastiRecursiveInterconnect_io_slaves_0_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = NastiRecursiveInterconnect_io_slaves_0_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = NastiRecursiveInterconnect_io_slaves_0_aw_bits_size;
  assign io_slaves_1_aw_bits_len = NastiRecursiveInterconnect_io_slaves_0_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = NastiRecursiveInterconnect_io_slaves_0_aw_bits_addr;
  assign io_slaves_1_aw_valid = NastiRecursiveInterconnect_io_slaves_0_aw_valid;
  assign io_slaves_2_r_ready = NastiRecursiveInterconnect_io_slaves_1_r_ready;
  assign io_slaves_2_ar_bits_user = NastiRecursiveInterconnect_io_slaves_1_ar_bits_user;
  assign io_slaves_2_ar_bits_id = NastiRecursiveInterconnect_io_slaves_1_ar_bits_id;
  assign io_slaves_2_ar_bits_region = NastiRecursiveInterconnect_io_slaves_1_ar_bits_region;
  assign io_slaves_2_ar_bits_qos = NastiRecursiveInterconnect_io_slaves_1_ar_bits_qos;
  assign io_slaves_2_ar_bits_prot = NastiRecursiveInterconnect_io_slaves_1_ar_bits_prot;
  assign io_slaves_2_ar_bits_cache = NastiRecursiveInterconnect_io_slaves_1_ar_bits_cache;
  assign io_slaves_2_ar_bits_lock = NastiRecursiveInterconnect_io_slaves_1_ar_bits_lock;
  assign io_slaves_2_ar_bits_burst = NastiRecursiveInterconnect_io_slaves_1_ar_bits_burst;
  assign io_slaves_2_ar_bits_size = NastiRecursiveInterconnect_io_slaves_1_ar_bits_size;
  assign io_slaves_2_ar_bits_len = NastiRecursiveInterconnect_io_slaves_1_ar_bits_len;
  assign io_slaves_2_ar_bits_addr = NastiRecursiveInterconnect_io_slaves_1_ar_bits_addr;
  assign io_slaves_2_ar_valid = NastiRecursiveInterconnect_io_slaves_1_ar_valid;
  assign io_slaves_2_b_ready = NastiRecursiveInterconnect_io_slaves_1_b_ready;
  assign io_slaves_2_w_bits_user = NastiRecursiveInterconnect_io_slaves_1_w_bits_user;
  assign io_slaves_2_w_bits_strb = NastiRecursiveInterconnect_io_slaves_1_w_bits_strb;
  assign io_slaves_2_w_bits_last = NastiRecursiveInterconnect_io_slaves_1_w_bits_last;
  assign io_slaves_2_w_bits_data = NastiRecursiveInterconnect_io_slaves_1_w_bits_data;
  assign io_slaves_2_w_valid = NastiRecursiveInterconnect_io_slaves_1_w_valid;
  assign io_slaves_2_aw_bits_user = NastiRecursiveInterconnect_io_slaves_1_aw_bits_user;
  assign io_slaves_2_aw_bits_id = NastiRecursiveInterconnect_io_slaves_1_aw_bits_id;
  assign io_slaves_2_aw_bits_region = NastiRecursiveInterconnect_io_slaves_1_aw_bits_region;
  assign io_slaves_2_aw_bits_qos = NastiRecursiveInterconnect_io_slaves_1_aw_bits_qos;
  assign io_slaves_2_aw_bits_prot = NastiRecursiveInterconnect_io_slaves_1_aw_bits_prot;
  assign io_slaves_2_aw_bits_cache = NastiRecursiveInterconnect_io_slaves_1_aw_bits_cache;
  assign io_slaves_2_aw_bits_lock = NastiRecursiveInterconnect_io_slaves_1_aw_bits_lock;
  assign io_slaves_2_aw_bits_burst = NastiRecursiveInterconnect_io_slaves_1_aw_bits_burst;
  assign io_slaves_2_aw_bits_size = NastiRecursiveInterconnect_io_slaves_1_aw_bits_size;
  assign io_slaves_2_aw_bits_len = NastiRecursiveInterconnect_io_slaves_1_aw_bits_len;
  assign io_slaves_2_aw_bits_addr = NastiRecursiveInterconnect_io_slaves_1_aw_bits_addr;
  assign io_slaves_2_aw_valid = NastiRecursiveInterconnect_io_slaves_1_aw_valid;
  assign io_slaves_3_r_ready = xbar_io_slaves_2_r_ready;
  assign io_slaves_3_ar_bits_user = xbar_io_slaves_2_ar_bits_user;
  assign io_slaves_3_ar_bits_id = xbar_io_slaves_2_ar_bits_id;
  assign io_slaves_3_ar_bits_region = xbar_io_slaves_2_ar_bits_region;
  assign io_slaves_3_ar_bits_qos = xbar_io_slaves_2_ar_bits_qos;
  assign io_slaves_3_ar_bits_prot = xbar_io_slaves_2_ar_bits_prot;
  assign io_slaves_3_ar_bits_cache = xbar_io_slaves_2_ar_bits_cache;
  assign io_slaves_3_ar_bits_lock = xbar_io_slaves_2_ar_bits_lock;
  assign io_slaves_3_ar_bits_burst = xbar_io_slaves_2_ar_bits_burst;
  assign io_slaves_3_ar_bits_size = xbar_io_slaves_2_ar_bits_size;
  assign io_slaves_3_ar_bits_len = xbar_io_slaves_2_ar_bits_len;
  assign io_slaves_3_ar_bits_addr = xbar_io_slaves_2_ar_bits_addr;
  assign io_slaves_3_ar_valid = xbar_io_slaves_2_ar_valid;
  assign io_slaves_3_b_ready = xbar_io_slaves_2_b_ready;
  assign io_slaves_3_w_bits_user = xbar_io_slaves_2_w_bits_user;
  assign io_slaves_3_w_bits_strb = xbar_io_slaves_2_w_bits_strb;
  assign io_slaves_3_w_bits_last = xbar_io_slaves_2_w_bits_last;
  assign io_slaves_3_w_bits_data = xbar_io_slaves_2_w_bits_data;
  assign io_slaves_3_w_valid = xbar_io_slaves_2_w_valid;
  assign io_slaves_3_aw_bits_user = xbar_io_slaves_2_aw_bits_user;
  assign io_slaves_3_aw_bits_id = xbar_io_slaves_2_aw_bits_id;
  assign io_slaves_3_aw_bits_region = xbar_io_slaves_2_aw_bits_region;
  assign io_slaves_3_aw_bits_qos = xbar_io_slaves_2_aw_bits_qos;
  assign io_slaves_3_aw_bits_prot = xbar_io_slaves_2_aw_bits_prot;
  assign io_slaves_3_aw_bits_cache = xbar_io_slaves_2_aw_bits_cache;
  assign io_slaves_3_aw_bits_lock = xbar_io_slaves_2_aw_bits_lock;
  assign io_slaves_3_aw_bits_burst = xbar_io_slaves_2_aw_bits_burst;
  assign io_slaves_3_aw_bits_size = xbar_io_slaves_2_aw_bits_size;
  assign io_slaves_3_aw_bits_len = xbar_io_slaves_2_aw_bits_len;
  assign io_slaves_3_aw_bits_addr = xbar_io_slaves_2_aw_bits_addr;
  assign io_slaves_3_aw_valid = xbar_io_slaves_2_aw_valid;
  assign io_masters_0_r_bits_user = xbar_io_masters_0_r_bits_user;
  assign io_masters_0_r_bits_id = xbar_io_masters_0_r_bits_id;
  assign io_masters_0_r_bits_last = xbar_io_masters_0_r_bits_last;
  assign io_masters_0_r_bits_data = xbar_io_masters_0_r_bits_data;
  assign io_masters_0_r_bits_resp = xbar_io_masters_0_r_bits_resp;
  assign io_masters_0_r_valid = xbar_io_masters_0_r_valid;
  assign io_masters_0_ar_ready = xbar_io_masters_0_ar_ready;
  assign io_masters_0_b_bits_user = xbar_io_masters_0_b_bits_user;
  assign io_masters_0_b_bits_id = xbar_io_masters_0_b_bits_id;
  assign io_masters_0_b_bits_resp = xbar_io_masters_0_b_bits_resp;
  assign io_masters_0_b_valid = xbar_io_masters_0_b_valid;
  assign io_masters_0_w_ready = xbar_io_masters_0_w_ready;
  assign io_masters_0_aw_ready = xbar_io_masters_0_aw_ready;
  assign io_masters_1_r_bits_user = xbar_io_masters_1_r_bits_user;
  assign io_masters_1_r_bits_id = xbar_io_masters_1_r_bits_id;
  assign io_masters_1_r_bits_last = xbar_io_masters_1_r_bits_last;
  assign io_masters_1_r_bits_data = xbar_io_masters_1_r_bits_data;
  assign io_masters_1_r_bits_resp = xbar_io_masters_1_r_bits_resp;
  assign io_masters_1_r_valid = xbar_io_masters_1_r_valid;
  assign io_masters_1_ar_ready = xbar_io_masters_1_ar_ready;
  assign io_masters_1_b_bits_user = xbar_io_masters_1_b_bits_user;
  assign io_masters_1_b_bits_id = xbar_io_masters_1_b_bits_id;
  assign io_masters_1_b_bits_resp = xbar_io_masters_1_b_bits_resp;
  assign io_masters_1_b_valid = xbar_io_masters_1_b_valid;
  assign io_masters_1_w_ready = xbar_io_masters_1_w_ready;
  assign io_masters_1_aw_ready = xbar_io_masters_1_aw_ready;
  NastiCrossbar_0 xbar(.clk(clk), .reset(reset),
       .io_masters_1_aw_ready( xbar_io_masters_1_aw_ready ),
       .io_masters_1_aw_valid( io_masters_1_aw_valid ),
       .io_masters_1_aw_bits_addr( io_masters_1_aw_bits_addr ),
       .io_masters_1_aw_bits_len( io_masters_1_aw_bits_len ),
       .io_masters_1_aw_bits_size( io_masters_1_aw_bits_size ),
       .io_masters_1_aw_bits_burst( io_masters_1_aw_bits_burst ),
       .io_masters_1_aw_bits_lock( io_masters_1_aw_bits_lock ),
       .io_masters_1_aw_bits_cache( io_masters_1_aw_bits_cache ),
       .io_masters_1_aw_bits_prot( io_masters_1_aw_bits_prot ),
       .io_masters_1_aw_bits_qos( io_masters_1_aw_bits_qos ),
       .io_masters_1_aw_bits_region( io_masters_1_aw_bits_region ),
       .io_masters_1_aw_bits_id( io_masters_1_aw_bits_id ),
       .io_masters_1_aw_bits_user( io_masters_1_aw_bits_user ),
       .io_masters_1_w_ready( xbar_io_masters_1_w_ready ),
       .io_masters_1_w_valid( io_masters_1_w_valid ),
       .io_masters_1_w_bits_data( io_masters_1_w_bits_data ),
       .io_masters_1_w_bits_last( io_masters_1_w_bits_last ),
       .io_masters_1_w_bits_strb( io_masters_1_w_bits_strb ),
       .io_masters_1_w_bits_user( io_masters_1_w_bits_user ),
       .io_masters_1_b_ready( io_masters_1_b_ready ),
       .io_masters_1_b_valid( xbar_io_masters_1_b_valid ),
       .io_masters_1_b_bits_resp( xbar_io_masters_1_b_bits_resp ),
       .io_masters_1_b_bits_id( xbar_io_masters_1_b_bits_id ),
       .io_masters_1_b_bits_user( xbar_io_masters_1_b_bits_user ),
       .io_masters_1_ar_ready( xbar_io_masters_1_ar_ready ),
       .io_masters_1_ar_valid( io_masters_1_ar_valid ),
       .io_masters_1_ar_bits_addr( io_masters_1_ar_bits_addr ),
       .io_masters_1_ar_bits_len( io_masters_1_ar_bits_len ),
       .io_masters_1_ar_bits_size( io_masters_1_ar_bits_size ),
       .io_masters_1_ar_bits_burst( io_masters_1_ar_bits_burst ),
       .io_masters_1_ar_bits_lock( io_masters_1_ar_bits_lock ),
       .io_masters_1_ar_bits_cache( io_masters_1_ar_bits_cache ),
       .io_masters_1_ar_bits_prot( io_masters_1_ar_bits_prot ),
       .io_masters_1_ar_bits_qos( io_masters_1_ar_bits_qos ),
       .io_masters_1_ar_bits_region( io_masters_1_ar_bits_region ),
       .io_masters_1_ar_bits_id( io_masters_1_ar_bits_id ),
       .io_masters_1_ar_bits_user( io_masters_1_ar_bits_user ),
       .io_masters_1_r_ready( io_masters_1_r_ready ),
       .io_masters_1_r_valid( xbar_io_masters_1_r_valid ),
       .io_masters_1_r_bits_resp( xbar_io_masters_1_r_bits_resp ),
       .io_masters_1_r_bits_data( xbar_io_masters_1_r_bits_data ),
       .io_masters_1_r_bits_last( xbar_io_masters_1_r_bits_last ),
       .io_masters_1_r_bits_id( xbar_io_masters_1_r_bits_id ),
       .io_masters_1_r_bits_user( xbar_io_masters_1_r_bits_user ),
       .io_masters_0_aw_ready( xbar_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( io_masters_0_aw_valid ),
       .io_masters_0_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_masters_0_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_masters_0_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_masters_0_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_masters_0_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_masters_0_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_masters_0_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_masters_0_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_masters_0_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_masters_0_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_masters_0_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_masters_0_w_ready( xbar_io_masters_0_w_ready ),
       .io_masters_0_w_valid( io_masters_0_w_valid ),
       .io_masters_0_w_bits_data( io_masters_0_w_bits_data ),
       .io_masters_0_w_bits_last( io_masters_0_w_bits_last ),
       .io_masters_0_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_masters_0_w_bits_user( io_masters_0_w_bits_user ),
       .io_masters_0_b_ready( io_masters_0_b_ready ),
       .io_masters_0_b_valid( xbar_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( xbar_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( xbar_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( xbar_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( xbar_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( io_masters_0_ar_valid ),
       .io_masters_0_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_masters_0_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_masters_0_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_masters_0_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_masters_0_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_masters_0_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_masters_0_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_masters_0_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_masters_0_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_masters_0_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_masters_0_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_masters_0_r_ready( io_masters_0_r_ready ),
       .io_masters_0_r_valid( xbar_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( xbar_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( xbar_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( xbar_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( xbar_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( xbar_io_masters_0_r_bits_user ),
       .io_slaves_2_aw_ready( io_slaves_3_aw_ready ),
       .io_slaves_2_aw_valid( xbar_io_slaves_2_aw_valid ),
       .io_slaves_2_aw_bits_addr( xbar_io_slaves_2_aw_bits_addr ),
       .io_slaves_2_aw_bits_len( xbar_io_slaves_2_aw_bits_len ),
       .io_slaves_2_aw_bits_size( xbar_io_slaves_2_aw_bits_size ),
       .io_slaves_2_aw_bits_burst( xbar_io_slaves_2_aw_bits_burst ),
       .io_slaves_2_aw_bits_lock( xbar_io_slaves_2_aw_bits_lock ),
       .io_slaves_2_aw_bits_cache( xbar_io_slaves_2_aw_bits_cache ),
       .io_slaves_2_aw_bits_prot( xbar_io_slaves_2_aw_bits_prot ),
       .io_slaves_2_aw_bits_qos( xbar_io_slaves_2_aw_bits_qos ),
       .io_slaves_2_aw_bits_region( xbar_io_slaves_2_aw_bits_region ),
       .io_slaves_2_aw_bits_id( xbar_io_slaves_2_aw_bits_id ),
       .io_slaves_2_aw_bits_user( xbar_io_slaves_2_aw_bits_user ),
       .io_slaves_2_w_ready( io_slaves_3_w_ready ),
       .io_slaves_2_w_valid( xbar_io_slaves_2_w_valid ),
       .io_slaves_2_w_bits_data( xbar_io_slaves_2_w_bits_data ),
       .io_slaves_2_w_bits_last( xbar_io_slaves_2_w_bits_last ),
       .io_slaves_2_w_bits_strb( xbar_io_slaves_2_w_bits_strb ),
       .io_slaves_2_w_bits_user( xbar_io_slaves_2_w_bits_user ),
       .io_slaves_2_b_ready( xbar_io_slaves_2_b_ready ),
       .io_slaves_2_b_valid( io_slaves_3_b_valid ),
       .io_slaves_2_b_bits_resp( io_slaves_3_b_bits_resp ),
       .io_slaves_2_b_bits_id( io_slaves_3_b_bits_id ),
       .io_slaves_2_b_bits_user( io_slaves_3_b_bits_user ),
       .io_slaves_2_ar_ready( io_slaves_3_ar_ready ),
       .io_slaves_2_ar_valid( xbar_io_slaves_2_ar_valid ),
       .io_slaves_2_ar_bits_addr( xbar_io_slaves_2_ar_bits_addr ),
       .io_slaves_2_ar_bits_len( xbar_io_slaves_2_ar_bits_len ),
       .io_slaves_2_ar_bits_size( xbar_io_slaves_2_ar_bits_size ),
       .io_slaves_2_ar_bits_burst( xbar_io_slaves_2_ar_bits_burst ),
       .io_slaves_2_ar_bits_lock( xbar_io_slaves_2_ar_bits_lock ),
       .io_slaves_2_ar_bits_cache( xbar_io_slaves_2_ar_bits_cache ),
       .io_slaves_2_ar_bits_prot( xbar_io_slaves_2_ar_bits_prot ),
       .io_slaves_2_ar_bits_qos( xbar_io_slaves_2_ar_bits_qos ),
       .io_slaves_2_ar_bits_region( xbar_io_slaves_2_ar_bits_region ),
       .io_slaves_2_ar_bits_id( xbar_io_slaves_2_ar_bits_id ),
       .io_slaves_2_ar_bits_user( xbar_io_slaves_2_ar_bits_user ),
       .io_slaves_2_r_ready( xbar_io_slaves_2_r_ready ),
       .io_slaves_2_r_valid( io_slaves_3_r_valid ),
       .io_slaves_2_r_bits_resp( io_slaves_3_r_bits_resp ),
       .io_slaves_2_r_bits_data( io_slaves_3_r_bits_data ),
       .io_slaves_2_r_bits_last( io_slaves_3_r_bits_last ),
       .io_slaves_2_r_bits_id( io_slaves_3_r_bits_id ),
       .io_slaves_2_r_bits_user( io_slaves_3_r_bits_user ),
       .io_slaves_1_aw_ready( NastiRecursiveInterconnect_io_masters_0_aw_ready ),
       .io_slaves_1_aw_valid( xbar_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( xbar_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( xbar_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( xbar_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( xbar_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( xbar_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( xbar_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( xbar_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( xbar_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( xbar_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( xbar_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( xbar_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( NastiRecursiveInterconnect_io_masters_0_w_ready ),
       .io_slaves_1_w_valid( xbar_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( xbar_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( xbar_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( xbar_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( xbar_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( xbar_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( NastiRecursiveInterconnect_io_masters_0_b_valid ),
       .io_slaves_1_b_bits_resp( NastiRecursiveInterconnect_io_masters_0_b_bits_resp ),
       .io_slaves_1_b_bits_id( NastiRecursiveInterconnect_io_masters_0_b_bits_id ),
       .io_slaves_1_b_bits_user( NastiRecursiveInterconnect_io_masters_0_b_bits_user ),
       .io_slaves_1_ar_ready( NastiRecursiveInterconnect_io_masters_0_ar_ready ),
       .io_slaves_1_ar_valid( xbar_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( xbar_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( xbar_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( xbar_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( xbar_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( xbar_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( xbar_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( xbar_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( xbar_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( xbar_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( xbar_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( xbar_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( xbar_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( NastiRecursiveInterconnect_io_masters_0_r_valid ),
       .io_slaves_1_r_bits_resp( NastiRecursiveInterconnect_io_masters_0_r_bits_resp ),
       .io_slaves_1_r_bits_data( NastiRecursiveInterconnect_io_masters_0_r_bits_data ),
       .io_slaves_1_r_bits_last( NastiRecursiveInterconnect_io_masters_0_r_bits_last ),
       .io_slaves_1_r_bits_id( NastiRecursiveInterconnect_io_masters_0_r_bits_id ),
       .io_slaves_1_r_bits_user( NastiRecursiveInterconnect_io_masters_0_r_bits_user ),
       .io_slaves_0_aw_ready( NastiMultiChannelRouter_io_master_aw_ready ),
       .io_slaves_0_aw_valid( xbar_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( xbar_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( xbar_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( xbar_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( xbar_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( xbar_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( xbar_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( xbar_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( xbar_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( xbar_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( xbar_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( xbar_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( NastiMultiChannelRouter_io_master_w_ready ),
       .io_slaves_0_w_valid( xbar_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( xbar_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( xbar_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( xbar_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( xbar_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( xbar_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( NastiMultiChannelRouter_io_master_b_valid ),
       .io_slaves_0_b_bits_resp( NastiMultiChannelRouter_io_master_b_bits_resp ),
       .io_slaves_0_b_bits_id( NastiMultiChannelRouter_io_master_b_bits_id ),
       .io_slaves_0_b_bits_user( NastiMultiChannelRouter_io_master_b_bits_user ),
       .io_slaves_0_ar_ready( NastiMultiChannelRouter_io_master_ar_ready ),
       .io_slaves_0_ar_valid( xbar_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( xbar_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( xbar_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( xbar_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( xbar_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( xbar_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( xbar_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( xbar_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( xbar_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( xbar_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( xbar_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( xbar_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( xbar_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( NastiMultiChannelRouter_io_master_r_valid ),
       .io_slaves_0_r_bits_resp( NastiMultiChannelRouter_io_master_r_bits_resp ),
       .io_slaves_0_r_bits_data( NastiMultiChannelRouter_io_master_r_bits_data ),
       .io_slaves_0_r_bits_last( NastiMultiChannelRouter_io_master_r_bits_last ),
       .io_slaves_0_r_bits_id( NastiMultiChannelRouter_io_master_r_bits_id ),
       .io_slaves_0_r_bits_user( NastiMultiChannelRouter_io_master_r_bits_user )
  );
  NastiMultiChannelRouter NastiMultiChannelRouter(
       .io_master_aw_ready( NastiMultiChannelRouter_io_master_aw_ready ),
       .io_master_aw_valid( xbar_io_slaves_0_aw_valid ),
       .io_master_aw_bits_addr( xbar_io_slaves_0_aw_bits_addr ),
       .io_master_aw_bits_len( xbar_io_slaves_0_aw_bits_len ),
       .io_master_aw_bits_size( xbar_io_slaves_0_aw_bits_size ),
       .io_master_aw_bits_burst( xbar_io_slaves_0_aw_bits_burst ),
       .io_master_aw_bits_lock( xbar_io_slaves_0_aw_bits_lock ),
       .io_master_aw_bits_cache( xbar_io_slaves_0_aw_bits_cache ),
       .io_master_aw_bits_prot( xbar_io_slaves_0_aw_bits_prot ),
       .io_master_aw_bits_qos( xbar_io_slaves_0_aw_bits_qos ),
       .io_master_aw_bits_region( xbar_io_slaves_0_aw_bits_region ),
       .io_master_aw_bits_id( xbar_io_slaves_0_aw_bits_id ),
       .io_master_aw_bits_user( xbar_io_slaves_0_aw_bits_user ),
       .io_master_w_ready( NastiMultiChannelRouter_io_master_w_ready ),
       .io_master_w_valid( xbar_io_slaves_0_w_valid ),
       .io_master_w_bits_data( xbar_io_slaves_0_w_bits_data ),
       .io_master_w_bits_last( xbar_io_slaves_0_w_bits_last ),
       .io_master_w_bits_strb( xbar_io_slaves_0_w_bits_strb ),
       .io_master_w_bits_user( xbar_io_slaves_0_w_bits_user ),
       .io_master_b_ready( xbar_io_slaves_0_b_ready ),
       .io_master_b_valid( NastiMultiChannelRouter_io_master_b_valid ),
       .io_master_b_bits_resp( NastiMultiChannelRouter_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiMultiChannelRouter_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiMultiChannelRouter_io_master_b_bits_user ),
       .io_master_ar_ready( NastiMultiChannelRouter_io_master_ar_ready ),
       .io_master_ar_valid( xbar_io_slaves_0_ar_valid ),
       .io_master_ar_bits_addr( xbar_io_slaves_0_ar_bits_addr ),
       .io_master_ar_bits_len( xbar_io_slaves_0_ar_bits_len ),
       .io_master_ar_bits_size( xbar_io_slaves_0_ar_bits_size ),
       .io_master_ar_bits_burst( xbar_io_slaves_0_ar_bits_burst ),
       .io_master_ar_bits_lock( xbar_io_slaves_0_ar_bits_lock ),
       .io_master_ar_bits_cache( xbar_io_slaves_0_ar_bits_cache ),
       .io_master_ar_bits_prot( xbar_io_slaves_0_ar_bits_prot ),
       .io_master_ar_bits_qos( xbar_io_slaves_0_ar_bits_qos ),
       .io_master_ar_bits_region( xbar_io_slaves_0_ar_bits_region ),
       .io_master_ar_bits_id( xbar_io_slaves_0_ar_bits_id ),
       .io_master_ar_bits_user( xbar_io_slaves_0_ar_bits_user ),
       .io_master_r_ready( xbar_io_slaves_0_r_ready ),
       .io_master_r_valid( NastiMultiChannelRouter_io_master_r_valid ),
       .io_master_r_bits_resp( NastiMultiChannelRouter_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiMultiChannelRouter_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiMultiChannelRouter_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiMultiChannelRouter_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiMultiChannelRouter_io_master_r_bits_user ),
       .io_slaves_0_aw_ready( io_slaves_0_aw_ready ),
       .io_slaves_0_aw_valid( NastiMultiChannelRouter_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( NastiMultiChannelRouter_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( NastiMultiChannelRouter_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( NastiMultiChannelRouter_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( NastiMultiChannelRouter_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( NastiMultiChannelRouter_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( NastiMultiChannelRouter_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( NastiMultiChannelRouter_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( NastiMultiChannelRouter_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( NastiMultiChannelRouter_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( NastiMultiChannelRouter_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( NastiMultiChannelRouter_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_slaves_0_w_ready ),
       .io_slaves_0_w_valid( NastiMultiChannelRouter_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( NastiMultiChannelRouter_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( NastiMultiChannelRouter_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( NastiMultiChannelRouter_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( NastiMultiChannelRouter_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( NastiMultiChannelRouter_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_slaves_0_b_valid ),
       .io_slaves_0_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slaves_0_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slaves_0_ar_ready( io_slaves_0_ar_ready ),
       .io_slaves_0_ar_valid( NastiMultiChannelRouter_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( NastiMultiChannelRouter_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( NastiMultiChannelRouter_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( NastiMultiChannelRouter_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( NastiMultiChannelRouter_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( NastiMultiChannelRouter_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( NastiMultiChannelRouter_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( NastiMultiChannelRouter_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( NastiMultiChannelRouter_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( NastiMultiChannelRouter_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( NastiMultiChannelRouter_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( NastiMultiChannelRouter_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( NastiMultiChannelRouter_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_slaves_0_r_valid ),
       .io_slaves_0_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slaves_0_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slaves_0_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slaves_0_r_bits_user( io_slaves_0_r_bits_user )
  );
  NastiRecursiveInterconnect NastiRecursiveInterconnect(.clk(clk), .reset(reset),
       .io_masters_0_aw_ready( NastiRecursiveInterconnect_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( xbar_io_slaves_1_aw_valid ),
       .io_masters_0_aw_bits_addr( xbar_io_slaves_1_aw_bits_addr ),
       .io_masters_0_aw_bits_len( xbar_io_slaves_1_aw_bits_len ),
       .io_masters_0_aw_bits_size( xbar_io_slaves_1_aw_bits_size ),
       .io_masters_0_aw_bits_burst( xbar_io_slaves_1_aw_bits_burst ),
       .io_masters_0_aw_bits_lock( xbar_io_slaves_1_aw_bits_lock ),
       .io_masters_0_aw_bits_cache( xbar_io_slaves_1_aw_bits_cache ),
       .io_masters_0_aw_bits_prot( xbar_io_slaves_1_aw_bits_prot ),
       .io_masters_0_aw_bits_qos( xbar_io_slaves_1_aw_bits_qos ),
       .io_masters_0_aw_bits_region( xbar_io_slaves_1_aw_bits_region ),
       .io_masters_0_aw_bits_id( xbar_io_slaves_1_aw_bits_id ),
       .io_masters_0_aw_bits_user( xbar_io_slaves_1_aw_bits_user ),
       .io_masters_0_w_ready( NastiRecursiveInterconnect_io_masters_0_w_ready ),
       .io_masters_0_w_valid( xbar_io_slaves_1_w_valid ),
       .io_masters_0_w_bits_data( xbar_io_slaves_1_w_bits_data ),
       .io_masters_0_w_bits_last( xbar_io_slaves_1_w_bits_last ),
       .io_masters_0_w_bits_strb( xbar_io_slaves_1_w_bits_strb ),
       .io_masters_0_w_bits_user( xbar_io_slaves_1_w_bits_user ),
       .io_masters_0_b_ready( xbar_io_slaves_1_b_ready ),
       .io_masters_0_b_valid( NastiRecursiveInterconnect_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( NastiRecursiveInterconnect_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( NastiRecursiveInterconnect_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( NastiRecursiveInterconnect_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( NastiRecursiveInterconnect_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( xbar_io_slaves_1_ar_valid ),
       .io_masters_0_ar_bits_addr( xbar_io_slaves_1_ar_bits_addr ),
       .io_masters_0_ar_bits_len( xbar_io_slaves_1_ar_bits_len ),
       .io_masters_0_ar_bits_size( xbar_io_slaves_1_ar_bits_size ),
       .io_masters_0_ar_bits_burst( xbar_io_slaves_1_ar_bits_burst ),
       .io_masters_0_ar_bits_lock( xbar_io_slaves_1_ar_bits_lock ),
       .io_masters_0_ar_bits_cache( xbar_io_slaves_1_ar_bits_cache ),
       .io_masters_0_ar_bits_prot( xbar_io_slaves_1_ar_bits_prot ),
       .io_masters_0_ar_bits_qos( xbar_io_slaves_1_ar_bits_qos ),
       .io_masters_0_ar_bits_region( xbar_io_slaves_1_ar_bits_region ),
       .io_masters_0_ar_bits_id( xbar_io_slaves_1_ar_bits_id ),
       .io_masters_0_ar_bits_user( xbar_io_slaves_1_ar_bits_user ),
       .io_masters_0_r_ready( xbar_io_slaves_1_r_ready ),
       .io_masters_0_r_valid( NastiRecursiveInterconnect_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( NastiRecursiveInterconnect_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( NastiRecursiveInterconnect_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( NastiRecursiveInterconnect_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( NastiRecursiveInterconnect_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( NastiRecursiveInterconnect_io_masters_0_r_bits_user ),
       .io_slaves_1_aw_ready( io_slaves_2_aw_ready ),
       .io_slaves_1_aw_valid( NastiRecursiveInterconnect_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( NastiRecursiveInterconnect_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( NastiRecursiveInterconnect_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( NastiRecursiveInterconnect_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( NastiRecursiveInterconnect_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( NastiRecursiveInterconnect_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( NastiRecursiveInterconnect_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( NastiRecursiveInterconnect_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( NastiRecursiveInterconnect_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( NastiRecursiveInterconnect_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( NastiRecursiveInterconnect_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( NastiRecursiveInterconnect_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( io_slaves_2_w_ready ),
       .io_slaves_1_w_valid( NastiRecursiveInterconnect_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( NastiRecursiveInterconnect_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( NastiRecursiveInterconnect_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( NastiRecursiveInterconnect_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( NastiRecursiveInterconnect_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( NastiRecursiveInterconnect_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( io_slaves_2_b_valid ),
       .io_slaves_1_b_bits_resp( io_slaves_2_b_bits_resp ),
       .io_slaves_1_b_bits_id( io_slaves_2_b_bits_id ),
       .io_slaves_1_b_bits_user( io_slaves_2_b_bits_user ),
       .io_slaves_1_ar_ready( io_slaves_2_ar_ready ),
       .io_slaves_1_ar_valid( NastiRecursiveInterconnect_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( NastiRecursiveInterconnect_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( NastiRecursiveInterconnect_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( NastiRecursiveInterconnect_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( NastiRecursiveInterconnect_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( NastiRecursiveInterconnect_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( NastiRecursiveInterconnect_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( NastiRecursiveInterconnect_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( NastiRecursiveInterconnect_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( NastiRecursiveInterconnect_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( NastiRecursiveInterconnect_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( NastiRecursiveInterconnect_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( NastiRecursiveInterconnect_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( io_slaves_2_r_valid ),
       .io_slaves_1_r_bits_resp( io_slaves_2_r_bits_resp ),
       .io_slaves_1_r_bits_data( io_slaves_2_r_bits_data ),
       .io_slaves_1_r_bits_last( io_slaves_2_r_bits_last ),
       .io_slaves_1_r_bits_id( io_slaves_2_r_bits_id ),
       .io_slaves_1_r_bits_user( io_slaves_2_r_bits_user ),
       .io_slaves_0_aw_ready( io_slaves_1_aw_ready ),
       .io_slaves_0_aw_valid( NastiRecursiveInterconnect_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( NastiRecursiveInterconnect_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( NastiRecursiveInterconnect_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( NastiRecursiveInterconnect_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( NastiRecursiveInterconnect_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( NastiRecursiveInterconnect_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( NastiRecursiveInterconnect_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( NastiRecursiveInterconnect_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( NastiRecursiveInterconnect_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( NastiRecursiveInterconnect_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( NastiRecursiveInterconnect_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( NastiRecursiveInterconnect_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_slaves_1_w_ready ),
       .io_slaves_0_w_valid( NastiRecursiveInterconnect_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( NastiRecursiveInterconnect_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( NastiRecursiveInterconnect_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( NastiRecursiveInterconnect_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( NastiRecursiveInterconnect_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( NastiRecursiveInterconnect_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_slaves_1_b_valid ),
       .io_slaves_0_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slaves_0_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slaves_0_ar_ready( io_slaves_1_ar_ready ),
       .io_slaves_0_ar_valid( NastiRecursiveInterconnect_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( NastiRecursiveInterconnect_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( NastiRecursiveInterconnect_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( NastiRecursiveInterconnect_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( NastiRecursiveInterconnect_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( NastiRecursiveInterconnect_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( NastiRecursiveInterconnect_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( NastiRecursiveInterconnect_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( NastiRecursiveInterconnect_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( NastiRecursiveInterconnect_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( NastiRecursiveInterconnect_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( NastiRecursiveInterconnect_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( NastiRecursiveInterconnect_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_slaves_1_r_valid ),
       .io_slaves_0_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slaves_0_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slaves_0_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slaves_0_r_bits_user( io_slaves_1_r_bits_user )
  );
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [3:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [3:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[3:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  wire T1;
  wire T2;
  wire T3;
  reg  last_grant;
  wire T52;
  wire T4;
  wire T5;
  reg  lockIdx;
  wire T53;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  reg  locked;
  wire T54;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  reg [1:0] R20;
  wire[1:0] T55;
  wire[1:0] T21;
  wire[127:0] T22;
  wire T23;
  wire[16:0] T24;
  wire[2:0] T25;
  wire T26;
  wire[1:0] T27;
  wire[3:0] T28;
  wire[25:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R20 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T2 ? 1'h1 : T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign T2 = io_in_1_valid & T3;
  assign T3 = last_grant < 1'h1;
  assign T52 = reset ? 1'h0 : T4;
  assign T4 = T5 ? chosen : last_grant;
  assign T5 = io_out_ready & io_out_valid;
  assign T53 = reset ? 1'h1 : T6;
  assign T6 = T9 ? T7 : lockIdx;
  assign T7 = T8 == 1'h0;
  assign T8 = io_in_0_ready & io_in_0_valid;
  assign T9 = T11 & T10;
  assign T10 = locked ^ 1'h1;
  assign T11 = T14 & T12;
  assign T12 = io_out_bits_is_builtin_type & T13;
  assign T13 = 3'h3 == io_out_bits_a_type;
  assign T14 = io_out_ready & io_out_valid;
  assign T54 = reset ? 1'h0 : T15;
  assign T15 = T17 ? 1'h0 : T16;
  assign T16 = T9 ? 1'h1 : locked;
  assign T17 = T14 & T18;
  assign T18 = T19 == 2'h0;
  assign T19 = R20 + 2'h1;
  assign T55 = reset ? 2'h0 : T21;
  assign T21 = T11 ? T19 : R20;
  assign io_out_bits_data = T22;
  assign T22 = T23 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T23 = chosen;
  assign io_out_bits_union = T24;
  assign T24 = T23 ? io_in_1_bits_union : io_in_0_bits_union;
  assign io_out_bits_a_type = T25;
  assign T25 = T23 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_is_builtin_type = T26;
  assign T26 = T23 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign io_out_bits_addr_beat = T27;
  assign T27 = T23 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_bits_client_xact_id = T28;
  assign T28 = T23 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T29;
  assign T29 = T23 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_valid = T30;
  assign T30 = T23 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = locked ? T41 : T33;
  assign T33 = T40 | T34;
  assign T34 = T35 ^ 1'h1;
  assign T35 = T38 | T36;
  assign T36 = io_in_1_valid & T37;
  assign T37 = last_grant < 1'h1;
  assign T38 = io_in_0_valid & T39;
  assign T39 = last_grant < 1'h0;
  assign T40 = last_grant < 1'h0;
  assign T41 = lockIdx == 1'h0;
  assign io_in_1_ready = T42;
  assign T42 = T43 & io_out_ready;
  assign T43 = locked ? T51 : T44;
  assign T44 = T48 | T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T47 | io_in_0_valid;
  assign T47 = T38 | T36;
  assign T48 = T50 & T49;
  assign T49 = last_grant < 1'h1;
  assign T50 = T38 ^ 1'h1;
  assign T51 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T5) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T9) begin
      lockIdx <= T7;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T17) begin
      locked <= 1'h0;
    end else if(T9) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R20 <= 2'h0;
    end else if(T11) begin
      R20 <= T19;
    end
  end
endmodule

module ReorderQueue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_data,
    input [3:0] io_enq_bits_tag,
    input  io_deq_valid,
    input [3:0] io_deq_tag,
    output io_deq_data,
    output io_deq_matches
);

  wire T0;
  wire roq_matches_8;
  wire T1;
  reg  roq_free_8;
  wire T182;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[15:0] T6;
  wire[3:0] T7;
  wire[3:0] roq_enq_addr;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  reg  roq_free_7;
  wire T183;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[15:0] T21;
  wire[3:0] T22;
  wire[3:0] roq_deq_addr;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  wire roq_matches_7;
  wire T30;
  wire T31;
  reg [3:0] roq_tags_7;
  wire[3:0] T32;
  wire T33;
  wire T34;
  wire[15:0] T35;
  wire[3:0] T36;
  wire roq_matches_6;
  wire T37;
  wire T38;
  reg [3:0] roq_tags_6;
  wire[3:0] T39;
  wire T40;
  wire T41;
  wire roq_matches_5;
  wire T42;
  wire T43;
  reg [3:0] roq_tags_5;
  wire[3:0] T44;
  wire T45;
  wire T46;
  wire roq_matches_4;
  wire T47;
  wire T48;
  reg [3:0] roq_tags_4;
  wire[3:0] T49;
  wire T50;
  wire T51;
  wire roq_matches_3;
  wire T52;
  wire T53;
  reg [3:0] roq_tags_3;
  wire[3:0] T54;
  wire T55;
  wire T56;
  wire roq_matches_2;
  wire T57;
  wire T58;
  reg [3:0] roq_tags_2;
  wire[3:0] T59;
  wire T60;
  wire T61;
  wire roq_matches_1;
  wire T62;
  wire T63;
  reg [3:0] roq_tags_1;
  wire[3:0] T64;
  wire T65;
  wire T66;
  wire roq_matches_0;
  wire T67;
  wire T68;
  reg [3:0] roq_tags_0;
  wire[3:0] T69;
  wire T70;
  wire T71;
  reg  roq_free_6;
  wire T184;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg  roq_free_5;
  wire T185;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  reg  roq_free_4;
  wire T186;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg  roq_free_3;
  wire T187;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  reg  roq_free_2;
  wire T188;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  reg  roq_free_1;
  wire T189;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg  roq_free_0;
  wire T190;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  reg [3:0] roq_tags_8;
  wire[3:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg  roq_data_0;
  wire T132;
  wire T133;
  wire T134;
  wire[15:0] T135;
  wire[3:0] T136;
  reg  roq_data_1;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire[3:0] T141;
  wire T142;
  reg  roq_data_2;
  wire T143;
  wire T144;
  wire T145;
  reg  roq_data_3;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg  roq_data_4;
  wire T153;
  wire T154;
  wire T155;
  reg  roq_data_5;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  reg  roq_data_6;
  wire T161;
  wire T162;
  wire T163;
  reg  roq_data_7;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  reg  roq_data_8;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    roq_free_8 = {1{$random}};
    roq_free_7 = {1{$random}};
    roq_tags_7 = {1{$random}};
    roq_tags_6 = {1{$random}};
    roq_tags_5 = {1{$random}};
    roq_tags_4 = {1{$random}};
    roq_tags_3 = {1{$random}};
    roq_tags_2 = {1{$random}};
    roq_tags_1 = {1{$random}};
    roq_tags_0 = {1{$random}};
    roq_free_6 = {1{$random}};
    roq_free_5 = {1{$random}};
    roq_free_4 = {1{$random}};
    roq_free_3 = {1{$random}};
    roq_free_2 = {1{$random}};
    roq_free_1 = {1{$random}};
    roq_free_0 = {1{$random}};
    roq_tags_8 = {1{$random}};
    roq_data_0 = {1{$random}};
    roq_data_1 = {1{$random}};
    roq_data_2 = {1{$random}};
    roq_data_3 = {1{$random}};
    roq_data_4 = {1{$random}};
    roq_data_5 = {1{$random}};
    roq_data_6 = {1{$random}};
    roq_data_7 = {1{$random}};
    roq_data_8 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_deq_matches = T0;
  assign T0 = T121 | roq_matches_8;
  assign roq_matches_8 = T117 & T1;
  assign T1 = roq_free_8 ^ 1'h1;
  assign T182 = reset ? 1'h1 : T2;
  assign T2 = T115 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : roq_free_8;
  assign T4 = T114 & T5;
  assign T5 = T6[4'h8:4'h8];
  assign T6 = 1'h1 << T7;
  assign T7 = roq_enq_addr;
  assign roq_enq_addr = roq_free_0 ? 4'h0 : T8;
  assign T8 = roq_free_1 ? 4'h1 : T9;
  assign T9 = roq_free_2 ? 4'h2 : T10;
  assign T10 = roq_free_3 ? 4'h3 : T11;
  assign T11 = roq_free_4 ? 4'h4 : T12;
  assign T12 = roq_free_5 ? 4'h5 : T13;
  assign T13 = roq_free_6 ? 4'h6 : T14;
  assign T14 = roq_free_7 ? 4'h7 : 4'h8;
  assign T183 = reset ? 1'h1 : T15;
  assign T15 = T19 ? 1'h1 : T16;
  assign T16 = T17 ? 1'h0 : roq_free_7;
  assign T17 = T114 & T18;
  assign T18 = T6[3'h7:3'h7];
  assign T19 = io_deq_valid & T20;
  assign T20 = T21[3'h7:3'h7];
  assign T21 = 1'h1 << T22;
  assign T22 = roq_deq_addr;
  assign roq_deq_addr = roq_matches_0 ? 4'h0 : T23;
  assign T23 = roq_matches_1 ? 4'h1 : T24;
  assign T24 = roq_matches_2 ? 4'h2 : T25;
  assign T25 = roq_matches_3 ? 4'h3 : T26;
  assign T26 = roq_matches_4 ? 4'h4 : T27;
  assign T27 = roq_matches_5 ? 4'h5 : T28;
  assign T28 = roq_matches_6 ? 4'h6 : T29;
  assign T29 = roq_matches_7 ? 4'h7 : 4'h8;
  assign roq_matches_7 = T31 & T30;
  assign T30 = roq_free_7 ^ 1'h1;
  assign T31 = roq_tags_7 == io_deq_tag;
  assign T32 = T33 ? io_enq_bits_tag : roq_tags_7;
  assign T33 = T114 & T34;
  assign T34 = T35[3'h7:3'h7];
  assign T35 = 1'h1 << T36;
  assign T36 = roq_enq_addr;
  assign roq_matches_6 = T38 & T37;
  assign T37 = roq_free_6 ^ 1'h1;
  assign T38 = roq_tags_6 == io_deq_tag;
  assign T39 = T40 ? io_enq_bits_tag : roq_tags_6;
  assign T40 = T114 & T41;
  assign T41 = T35[3'h6:3'h6];
  assign roq_matches_5 = T43 & T42;
  assign T42 = roq_free_5 ^ 1'h1;
  assign T43 = roq_tags_5 == io_deq_tag;
  assign T44 = T45 ? io_enq_bits_tag : roq_tags_5;
  assign T45 = T114 & T46;
  assign T46 = T35[3'h5:3'h5];
  assign roq_matches_4 = T48 & T47;
  assign T47 = roq_free_4 ^ 1'h1;
  assign T48 = roq_tags_4 == io_deq_tag;
  assign T49 = T50 ? io_enq_bits_tag : roq_tags_4;
  assign T50 = T114 & T51;
  assign T51 = T35[3'h4:3'h4];
  assign roq_matches_3 = T53 & T52;
  assign T52 = roq_free_3 ^ 1'h1;
  assign T53 = roq_tags_3 == io_deq_tag;
  assign T54 = T55 ? io_enq_bits_tag : roq_tags_3;
  assign T55 = T114 & T56;
  assign T56 = T35[2'h3:2'h3];
  assign roq_matches_2 = T58 & T57;
  assign T57 = roq_free_2 ^ 1'h1;
  assign T58 = roq_tags_2 == io_deq_tag;
  assign T59 = T60 ? io_enq_bits_tag : roq_tags_2;
  assign T60 = T114 & T61;
  assign T61 = T35[2'h2:2'h2];
  assign roq_matches_1 = T63 & T62;
  assign T62 = roq_free_1 ^ 1'h1;
  assign T63 = roq_tags_1 == io_deq_tag;
  assign T64 = T65 ? io_enq_bits_tag : roq_tags_1;
  assign T65 = T114 & T66;
  assign T66 = T35[1'h1:1'h1];
  assign roq_matches_0 = T68 & T67;
  assign T67 = roq_free_0 ^ 1'h1;
  assign T68 = roq_tags_0 == io_deq_tag;
  assign T69 = T70 ? io_enq_bits_tag : roq_tags_0;
  assign T70 = T114 & T71;
  assign T71 = T35[1'h0:1'h0];
  assign T184 = reset ? 1'h1 : T72;
  assign T72 = T76 ? 1'h1 : T73;
  assign T73 = T74 ? 1'h0 : roq_free_6;
  assign T74 = T114 & T75;
  assign T75 = T6[3'h6:3'h6];
  assign T76 = io_deq_valid & T77;
  assign T77 = T21[3'h6:3'h6];
  assign T185 = reset ? 1'h1 : T78;
  assign T78 = T82 ? 1'h1 : T79;
  assign T79 = T80 ? 1'h0 : roq_free_5;
  assign T80 = T114 & T81;
  assign T81 = T6[3'h5:3'h5];
  assign T82 = io_deq_valid & T83;
  assign T83 = T21[3'h5:3'h5];
  assign T186 = reset ? 1'h1 : T84;
  assign T84 = T88 ? 1'h1 : T85;
  assign T85 = T86 ? 1'h0 : roq_free_4;
  assign T86 = T114 & T87;
  assign T87 = T6[3'h4:3'h4];
  assign T88 = io_deq_valid & T89;
  assign T89 = T21[3'h4:3'h4];
  assign T187 = reset ? 1'h1 : T90;
  assign T90 = T94 ? 1'h1 : T91;
  assign T91 = T92 ? 1'h0 : roq_free_3;
  assign T92 = T114 & T93;
  assign T93 = T6[2'h3:2'h3];
  assign T94 = io_deq_valid & T95;
  assign T95 = T21[2'h3:2'h3];
  assign T188 = reset ? 1'h1 : T96;
  assign T96 = T100 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : roq_free_2;
  assign T98 = T114 & T99;
  assign T99 = T6[2'h2:2'h2];
  assign T100 = io_deq_valid & T101;
  assign T101 = T21[2'h2:2'h2];
  assign T189 = reset ? 1'h1 : T102;
  assign T102 = T106 ? 1'h1 : T103;
  assign T103 = T104 ? 1'h0 : roq_free_1;
  assign T104 = T114 & T105;
  assign T105 = T6[1'h1:1'h1];
  assign T106 = io_deq_valid & T107;
  assign T107 = T21[1'h1:1'h1];
  assign T190 = reset ? 1'h1 : T108;
  assign T108 = T112 ? 1'h1 : T109;
  assign T109 = T110 ? 1'h0 : roq_free_0;
  assign T110 = T114 & T111;
  assign T111 = T6[1'h0:1'h0];
  assign T112 = io_deq_valid & T113;
  assign T113 = T21[1'h0:1'h0];
  assign T114 = io_enq_valid & io_enq_ready;
  assign T115 = io_deq_valid & T116;
  assign T116 = T21[4'h8:4'h8];
  assign T117 = roq_tags_8 == io_deq_tag;
  assign T118 = T119 ? io_enq_bits_tag : roq_tags_8;
  assign T119 = T114 & T120;
  assign T120 = T35[4'h8:4'h8];
  assign T121 = T122 | roq_matches_7;
  assign T122 = T123 | roq_matches_6;
  assign T123 = T124 | roq_matches_5;
  assign T124 = T125 | roq_matches_4;
  assign T125 = T126 | roq_matches_3;
  assign T126 = T127 | roq_matches_2;
  assign T127 = roq_matches_0 | roq_matches_1;
  assign io_deq_data = T128;
  assign T128 = T173 ? roq_data_8 : T129;
  assign T129 = T169 ? T151 : T130;
  assign T130 = T150 ? T142 : T131;
  assign T131 = T140 ? roq_data_1 : roq_data_0;
  assign T132 = T133 ? io_enq_bits_data : roq_data_0;
  assign T133 = T114 & T134;
  assign T134 = T135[1'h0:1'h0];
  assign T135 = 1'h1 << T136;
  assign T136 = roq_enq_addr;
  assign T137 = T138 ? io_enq_bits_data : roq_data_1;
  assign T138 = T114 & T139;
  assign T139 = T135[1'h1:1'h1];
  assign T140 = T141[1'h0:1'h0];
  assign T141 = roq_deq_addr;
  assign T142 = T149 ? roq_data_3 : roq_data_2;
  assign T143 = T144 ? io_enq_bits_data : roq_data_2;
  assign T144 = T114 & T145;
  assign T145 = T135[2'h2:2'h2];
  assign T146 = T147 ? io_enq_bits_data : roq_data_3;
  assign T147 = T114 & T148;
  assign T148 = T135[2'h3:2'h3];
  assign T149 = T141[1'h0:1'h0];
  assign T150 = T141[1'h1:1'h1];
  assign T151 = T168 ? T160 : T152;
  assign T152 = T159 ? roq_data_5 : roq_data_4;
  assign T153 = T154 ? io_enq_bits_data : roq_data_4;
  assign T154 = T114 & T155;
  assign T155 = T135[3'h4:3'h4];
  assign T156 = T157 ? io_enq_bits_data : roq_data_5;
  assign T157 = T114 & T158;
  assign T158 = T135[3'h5:3'h5];
  assign T159 = T141[1'h0:1'h0];
  assign T160 = T167 ? roq_data_7 : roq_data_6;
  assign T161 = T162 ? io_enq_bits_data : roq_data_6;
  assign T162 = T114 & T163;
  assign T163 = T135[3'h6:3'h6];
  assign T164 = T165 ? io_enq_bits_data : roq_data_7;
  assign T165 = T114 & T166;
  assign T166 = T135[3'h7:3'h7];
  assign T167 = T141[1'h0:1'h0];
  assign T168 = T141[1'h1:1'h1];
  assign T169 = T141[2'h2:2'h2];
  assign T170 = T171 ? io_enq_bits_data : roq_data_8;
  assign T171 = T114 & T172;
  assign T172 = T135[4'h8:4'h8];
  assign T173 = T141[2'h3:2'h3];
  assign io_enq_ready = T174;
  assign T174 = T175 | roq_free_8;
  assign T175 = T176 | roq_free_7;
  assign T176 = T177 | roq_free_6;
  assign T177 = T178 | roq_free_5;
  assign T178 = T179 | roq_free_4;
  assign T179 = T180 | roq_free_3;
  assign T180 = T181 | roq_free_2;
  assign T181 = roq_free_0 | roq_free_1;

  always @(posedge clk) begin
    if(reset) begin
      roq_free_8 <= 1'h1;
    end else if(T115) begin
      roq_free_8 <= 1'h1;
    end else if(T4) begin
      roq_free_8 <= 1'h0;
    end
    if(reset) begin
      roq_free_7 <= 1'h1;
    end else if(T19) begin
      roq_free_7 <= 1'h1;
    end else if(T17) begin
      roq_free_7 <= 1'h0;
    end
    if(T33) begin
      roq_tags_7 <= io_enq_bits_tag;
    end
    if(T40) begin
      roq_tags_6 <= io_enq_bits_tag;
    end
    if(T45) begin
      roq_tags_5 <= io_enq_bits_tag;
    end
    if(T50) begin
      roq_tags_4 <= io_enq_bits_tag;
    end
    if(T55) begin
      roq_tags_3 <= io_enq_bits_tag;
    end
    if(T60) begin
      roq_tags_2 <= io_enq_bits_tag;
    end
    if(T65) begin
      roq_tags_1 <= io_enq_bits_tag;
    end
    if(T70) begin
      roq_tags_0 <= io_enq_bits_tag;
    end
    if(reset) begin
      roq_free_6 <= 1'h1;
    end else if(T76) begin
      roq_free_6 <= 1'h1;
    end else if(T74) begin
      roq_free_6 <= 1'h0;
    end
    if(reset) begin
      roq_free_5 <= 1'h1;
    end else if(T82) begin
      roq_free_5 <= 1'h1;
    end else if(T80) begin
      roq_free_5 <= 1'h0;
    end
    if(reset) begin
      roq_free_4 <= 1'h1;
    end else if(T88) begin
      roq_free_4 <= 1'h1;
    end else if(T86) begin
      roq_free_4 <= 1'h0;
    end
    if(reset) begin
      roq_free_3 <= 1'h1;
    end else if(T94) begin
      roq_free_3 <= 1'h1;
    end else if(T92) begin
      roq_free_3 <= 1'h0;
    end
    if(reset) begin
      roq_free_2 <= 1'h1;
    end else if(T100) begin
      roq_free_2 <= 1'h1;
    end else if(T98) begin
      roq_free_2 <= 1'h0;
    end
    if(reset) begin
      roq_free_1 <= 1'h1;
    end else if(T106) begin
      roq_free_1 <= 1'h1;
    end else if(T104) begin
      roq_free_1 <= 1'h0;
    end
    if(reset) begin
      roq_free_0 <= 1'h1;
    end else if(T112) begin
      roq_free_0 <= 1'h1;
    end else if(T110) begin
      roq_free_0 <= 1'h0;
    end
    if(T119) begin
      roq_tags_8 <= io_enq_bits_tag;
    end
    if(T133) begin
      roq_data_0 <= io_enq_bits_data;
    end
    if(T138) begin
      roq_data_1 <= io_enq_bits_data;
    end
    if(T144) begin
      roq_data_2 <= io_enq_bits_data;
    end
    if(T147) begin
      roq_data_3 <= io_enq_bits_data;
    end
    if(T154) begin
      roq_data_4 <= io_enq_bits_data;
    end
    if(T157) begin
      roq_data_5 <= io_enq_bits_data;
    end
    if(T162) begin
      roq_data_6 <= io_enq_bits_data;
    end
    if(T165) begin
      roq_data_7 <= io_enq_bits_data;
    end
    if(T171) begin
      roq_data_8 <= io_enq_bits_data;
    end
  end
endmodule

module ClientTileLinkIOUnwrapper(input clk, input reset,
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [3:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[3:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_in_probe_ready,
    output io_in_probe_valid,
    //output[25:0] io_in_probe_bits_addr_block
    //output[1:0] io_in_probe_bits_p_type
    output io_in_release_ready,
    input  io_in_release_valid,
    input [1:0] io_in_release_bits_addr_beat,
    input [25:0] io_in_release_bits_addr_block,
    input [3:0] io_in_release_bits_client_xact_id,
    input [2:0] io_in_release_bits_r_type,
    input  io_in_release_bits_voluntary,
    input [127:0] io_in_release_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[3:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [3:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire rel_roq_enq;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire acq_roq_enq;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire[127:0] T31;
  wire[16:0] T32;
  wire[16:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire T36;
  wire[1:0] T37;
  wire[3:0] T38;
  wire[25:0] T39;
  wire T40;
  wire acq_roq_ready;
  wire T41;
  wire[127:0] T42;
  wire[16:0] T43;
  wire[16:0] T44;
  wire T45;
  wire[15:0] T46;
  wire[15:0] T47;
  wire[2:0] T48;
  wire T49;
  wire[1:0] T50;
  wire[3:0] T51;
  wire[25:0] T52;
  wire T53;
  wire rel_roq_ready;
  wire T54;
  wire T55;
  wire[127:0] T56;
  wire[127:0] rel_grant_data;
  wire[127:0] acq_grant_data;
  wire[3:0] T57;
  wire[3:0] rel_grant_g_type;
  wire[3:0] T58;
  wire[3:0] acq_grant_g_type;
  wire[3:0] T59;
  wire T60;
  wire rel_grant_is_builtin_type;
  wire acq_grant_is_builtin_type;
  wire T61;
  wire rel_grant_manager_xact_id;
  wire acq_grant_manager_xact_id;
  wire[3:0] T62;
  wire[3:0] rel_grant_client_xact_id;
  wire[3:0] acq_grant_client_xact_id;
  wire[1:0] T63;
  wire[1:0] rel_grant_addr_beat;
  wire[1:0] acq_grant_addr_beat;
  wire T64;
  wire acqArb_io_in_1_ready;
  wire acqArb_io_in_0_ready;
  wire acqArb_io_out_valid;
  wire[25:0] acqArb_io_out_bits_addr_block;
  wire[3:0] acqArb_io_out_bits_client_xact_id;
  wire[1:0] acqArb_io_out_bits_addr_beat;
  wire acqArb_io_out_bits_is_builtin_type;
  wire[2:0] acqArb_io_out_bits_a_type;
  wire[16:0] acqArb_io_out_bits_union;
  wire[127:0] acqArb_io_out_bits_data;
  wire acqRoq_io_enq_ready;
  wire acqRoq_io_deq_data;
  wire acqRoq_io_deq_matches;
  wire relRoq_io_enq_ready;
  wire relRoq_io_deq_data;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_in_probe_bits_p_type = {1{$random}};
//  assign io_in_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T7 & T1;
  assign T1 = T3 | T2;
  assign T2 = io_out_grant_bits_addr_beat == 2'h3;
  assign T3 = T4 ^ 1'h1;
  assign T4 = io_out_grant_bits_is_builtin_type ? T6 : T5;
  assign T5 = 4'h0 == io_out_grant_bits_g_type;
  assign T6 = 4'h5 == io_out_grant_bits_g_type;
  assign T7 = io_out_grant_ready & io_out_grant_valid;
  assign T8 = T16 & rel_roq_enq;
  assign rel_roq_enq = T10 | T9;
  assign T9 = io_in_release_bits_addr_beat == 2'h0;
  assign T10 = T11 ^ 1'h1;
  assign T11 = T13 | T12;
  assign T12 = 3'h2 == io_in_release_bits_r_type;
  assign T13 = T15 | T14;
  assign T14 = 3'h1 == io_in_release_bits_r_type;
  assign T15 = 3'h0 == io_in_release_bits_r_type;
  assign T16 = io_in_release_valid & acqArb_io_in_1_ready;
  assign T17 = T24 & T18;
  assign T18 = T20 | T19;
  assign T19 = io_out_grant_bits_addr_beat == 2'h3;
  assign T20 = T21 ^ 1'h1;
  assign T21 = io_out_grant_bits_is_builtin_type ? T23 : T22;
  assign T22 = 4'h0 == io_out_grant_bits_g_type;
  assign T23 = 4'h5 == io_out_grant_bits_g_type;
  assign T24 = io_out_grant_ready & io_out_grant_valid;
  assign T25 = T30 & acq_roq_enq;
  assign acq_roq_enq = T27 | T26;
  assign T26 = io_in_acquire_bits_addr_beat == 2'h0;
  assign T27 = T28 ^ 1'h1;
  assign T28 = io_in_acquire_bits_is_builtin_type & T29;
  assign T29 = 3'h3 == io_in_acquire_bits_a_type;
  assign T30 = io_in_acquire_valid & acqArb_io_in_0_ready;
  assign T31 = io_in_acquire_bits_data;
  assign T32 = T33;
  assign T33 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_union : 17'h1c1;
  assign T34 = T35;
  assign T35 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_a_type : 3'h1;
  assign T36 = 1'h1;
  assign T37 = io_in_acquire_bits_addr_beat;
  assign T38 = io_in_acquire_bits_client_xact_id;
  assign T39 = io_in_acquire_bits_addr_block;
  assign T40 = io_in_acquire_valid & acq_roq_ready;
  assign acq_roq_ready = T41 | acqRoq_io_enq_ready;
  assign T41 = acq_roq_enq ^ 1'h1;
  assign T42 = io_in_release_bits_data;
  assign T43 = T44;
  assign T44 = {T47, T45};
  assign T45 = T47 != T46;
  assign T46 = 16'hffff;
  assign T47 = 16'hffff;
  assign T48 = 3'h3;
  assign T49 = 1'h1;
  assign T50 = io_in_release_bits_addr_beat;
  assign T51 = io_in_release_bits_client_xact_id;
  assign T52 = io_in_release_bits_addr_block;
  assign T53 = io_in_release_valid & rel_roq_ready;
  assign rel_roq_ready = T54 | relRoq_io_enq_ready;
  assign T54 = rel_roq_enq ^ 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_data = acqArb_io_out_bits_data;
  assign io_out_acquire_bits_union = acqArb_io_out_bits_union;
  assign io_out_acquire_bits_a_type = acqArb_io_out_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = acqArb_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = acqArb_io_out_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = acqArb_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = acqArb_io_out_bits_addr_block;
  assign io_out_acquire_valid = acqArb_io_out_valid;
  assign io_in_release_ready = T55;
  assign T55 = rel_roq_ready & acqArb_io_in_1_ready;
  assign io_in_probe_valid = 1'h0;
  assign io_in_grant_bits_data = T56;
  assign T56 = acqRoq_io_deq_matches ? acq_grant_data : rel_grant_data;
  assign rel_grant_data = io_out_grant_bits_data;
  assign acq_grant_data = io_out_grant_bits_data;
  assign io_in_grant_bits_g_type = T57;
  assign T57 = acqRoq_io_deq_matches ? acq_grant_g_type : rel_grant_g_type;
  assign rel_grant_g_type = T58;
  assign T58 = relRoq_io_deq_data ? 4'h0 : io_out_grant_bits_g_type;
  assign acq_grant_g_type = T59;
  assign T59 = acqRoq_io_deq_data ? io_out_grant_bits_g_type : 4'h0;
  assign io_in_grant_bits_is_builtin_type = T60;
  assign T60 = acqRoq_io_deq_matches ? acq_grant_is_builtin_type : rel_grant_is_builtin_type;
  assign rel_grant_is_builtin_type = 1'h1;
  assign acq_grant_is_builtin_type = acqRoq_io_deq_data;
  assign io_in_grant_bits_manager_xact_id = T61;
  assign T61 = acqRoq_io_deq_matches ? acq_grant_manager_xact_id : rel_grant_manager_xact_id;
  assign rel_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign acq_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = T62;
  assign T62 = acqRoq_io_deq_matches ? acq_grant_client_xact_id : rel_grant_client_xact_id;
  assign rel_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign acq_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_addr_beat = T63;
  assign T63 = acqRoq_io_deq_matches ? acq_grant_addr_beat : rel_grant_addr_beat;
  assign rel_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign acq_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = T64;
  assign T64 = acq_roq_ready & acqArb_io_in_0_ready;
  LockingRRArbiter_4 acqArb(.clk(clk), .reset(reset),
       .io_in_1_ready( acqArb_io_in_1_ready ),
       .io_in_1_valid( T53 ),
       .io_in_1_bits_addr_block( T52 ),
       .io_in_1_bits_client_xact_id( T51 ),
       .io_in_1_bits_addr_beat( T50 ),
       .io_in_1_bits_is_builtin_type( T49 ),
       .io_in_1_bits_a_type( T48 ),
       .io_in_1_bits_union( T43 ),
       .io_in_1_bits_data( T42 ),
       .io_in_0_ready( acqArb_io_in_0_ready ),
       .io_in_0_valid( T40 ),
       .io_in_0_bits_addr_block( T39 ),
       .io_in_0_bits_client_xact_id( T38 ),
       .io_in_0_bits_addr_beat( T37 ),
       .io_in_0_bits_is_builtin_type( T36 ),
       .io_in_0_bits_a_type( T34 ),
       .io_in_0_bits_union( T32 ),
       .io_in_0_bits_data( T31 ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( acqArb_io_out_valid ),
       .io_out_bits_addr_block( acqArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( acqArb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( acqArb_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( acqArb_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( acqArb_io_out_bits_a_type ),
       .io_out_bits_union( acqArb_io_out_bits_union ),
       .io_out_bits_data( acqArb_io_out_bits_data )
       //.io_chosen(  )
  );
  ReorderQueue_0 acqRoq(.clk(clk), .reset(reset),
       .io_enq_ready( acqRoq_io_enq_ready ),
       .io_enq_valid( T25 ),
       .io_enq_bits_data( io_in_acquire_bits_is_builtin_type ),
       .io_enq_bits_tag( io_in_acquire_bits_client_xact_id ),
       .io_deq_valid( T17 ),
       .io_deq_tag( io_out_grant_bits_client_xact_id ),
       .io_deq_data( acqRoq_io_deq_data ),
       .io_deq_matches( acqRoq_io_deq_matches )
  );
  ReorderQueue_0 relRoq(.clk(clk), .reset(reset),
       .io_enq_ready( relRoq_io_enq_ready ),
       .io_enq_valid( T8 ),
       .io_enq_bits_data( io_in_release_bits_voluntary ),
       .io_enq_bits_tag( io_in_release_bits_client_xact_id ),
       .io_deq_valid( T0 ),
       .io_deq_tag( io_out_grant_bits_client_xact_id ),
       .io_deq_data( relRoq_io_deq_data )
       //.io_deq_matches(  )
  );
endmodule

module TileLinkIONarrower(input clk, input reset,
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [3:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[3:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[3:0] io_out_acquire_bits_client_xact_id,
    output[2:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[11:0] io_out_acquire_bits_union,
    output[63:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [2:0] io_out_grant_bits_addr_beat,
    input [3:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [63:0] io_out_grant_bits_data
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[2:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg[0:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire[7:0] T28;
  wire[15:0] T29;
  wire[15:0] T30;
  wire[15:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[15:0] T37;
  wire[15:0] T38;
  wire[7:0] T39;
  wire[7:0] T302;
  wire T40;
  wire[1:0] T41;
  wire T42;
  wire[3:0] T43;
  wire[7:0] T44;
  wire[7:0] T303;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire[15:0] T50;
  wire[15:0] T51;
  wire[15:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[15:0] T58;
  wire[15:0] T59;
  wire[7:0] T60;
  wire[7:0] T304;
  wire T61;
  wire[1:0] T62;
  wire T63;
  wire[3:0] T64;
  wire[7:0] T65;
  wire[7:0] T305;
  wire T66;
  wire T67;
  wire T68;
  wire[1:0] T306;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[31:0] T78;
  wire[5:0] T79;
  wire[3:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  reg  R89;
  wire T307;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  reg  R94;
  wire T308;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire[63:0] T309;
  wire[127:0] T101;
  wire[127:0] T102;
  wire[127:0] T103;
  wire[127:0] T104;
  wire[127:0] T310;
  wire[63:0] T105;
  wire[127:0] T311;
  wire[63:0] T106;
  wire[63:0] T107;
  wire[63:0] T108;
  wire[63:0] T109;
  wire T110;
  wire[63:0] T111;
  wire[63:0] T112;
  wire T113;
  wire[127:0] T312;
  wire[63:0] T114;
  wire T115;
  wire[127:0] T313;
  wire[63:0] T116;
  wire[63:0] T117;
  reg [127:0] R118;
  wire[127:0] T119;
  wire[127:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire[127:0] T314;
  wire[63:0] T124;
  wire T125;
  reg  R126;
  wire T315;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  reg  R131;
  wire T316;
  wire T132;
  wire T133;
  wire[11:0] T317;
  wire[16:0] T134;
  wire[16:0] T135;
  wire[16:0] T136;
  wire[16:0] T137;
  wire[16:0] T318;
  wire[11:0] T138;
  wire[11:0] T139;
  wire[5:0] T140;
  wire T141;
  wire[5:0] T142;
  wire[2:0] T143;
  wire[2:0] T144;
  wire[31:0] T145;
  wire[5:0] T146;
  wire[3:0] T147;
  wire[16:0] T319;
  wire[11:0] T148;
  wire[11:0] T320;
  wire[8:0] T149;
  wire[7:0] T150;
  wire[7:0] T151;
  wire T152;
  wire[7:0] T153;
  wire T154;
  wire[16:0] T321;
  wire[11:0] T155;
  wire[11:0] T322;
  wire[8:0] T156;
  wire[5:0] T157;
  wire T158;
  wire[16:0] T323;
  wire[11:0] T159;
  wire[11:0] T324;
  wire[8:0] T160;
  wire T161;
  wire[7:0] T162;
  wire[7:0] T163;
  reg [15:0] R164;
  wire[15:0] T165;
  wire[15:0] T166;
  wire[15:0] T167;
  wire[15:0] T168;
  wire[15:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire[15:0] T175;
  wire[15:0] T176;
  wire[7:0] T177;
  wire[7:0] T325;
  wire T178;
  wire[1:0] T179;
  wire T180;
  wire[3:0] T181;
  wire[7:0] T182;
  wire[7:0] T326;
  wire T183;
  wire T184;
  wire T185;
  wire[15:0] T327;
  wire[7:0] T186;
  wire[2:0] T187;
  wire[2:0] T188;
  wire[2:0] T189;
  wire[2:0] T190;
  wire[2:0] T191;
  wire[2:0] T192;
  wire[2:0] T193;
  wire[2:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire[2:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[2:0] T206;
  wire[2:0] T328;
  wire[2:0] T207;
  wire[2:0] T208;
  wire[31:0] T209;
  wire[5:0] T210;
  wire[3:0] T211;
  wire[2:0] T212;
  wire[2:0] T213;
  wire T329;
  wire T330;
  wire[2:0] T215;
  wire[2:0] T216;
  wire[2:0] T217;
  reg [1:0] R218;
  wire[1:0] T219;
  wire[3:0] T220;
  wire[3:0] T221;
  wire[3:0] T222;
  wire[3:0] T223;
  wire[3:0] T224;
  wire[3:0] T225;
  wire[3:0] T226;
  wire[3:0] T227;
  reg [3:0] R228;
  wire[3:0] T229;
  wire[25:0] T230;
  wire[25:0] T231;
  wire[25:0] T232;
  wire[25:0] T233;
  wire[25:0] T234;
  wire[25:0] T235;
  wire[25:0] T236;
  wire[25:0] T237;
  reg [25:0] R238;
  wire[25:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire[127:0] T247;
  wire[127:0] T248;
  wire[127:0] T331;
  wire[127:0] T249;
  wire[127:0] T332;
  wire[190:0] T250;
  wire[6:0] T251;
  wire[127:0] T252;
  wire[127:0] T253;
  wire[127:0] T254;
  reg [63:0] R255;
  wire[63:0] T256;
  wire T257;
  wire T258;
  wire[1:0] T259;
  wire T260;
  reg [63:0] R261;
  wire[63:0] T262;
  wire T263;
  wire T264;
  wire[3:0] T265;
  wire[3:0] T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  reg  R277;
  wire T278;
  wire[3:0] T279;
  wire[3:0] T280;
  wire[3:0] T281;
  wire[3:0] T282;
  reg [3:0] R283;
  wire[3:0] T284;
  wire[1:0] T333;
  wire[2:0] T285;
  wire[2:0] T286;
  wire[2:0] T334;
  wire[1:0] T287;
  wire[1:0] T335;
  wire[2:0] T336;
  wire[1:0] T288;
  reg [1:0] R289;
  wire[1:0] T337;
  wire[1:0] T290;
  wire[1:0] T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire ReorderQueue_io_enq_ready;
  wire ReorderQueue_io_deq_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T19 = 1'b0;
    R89 = {1{$random}};
    R94 = {1{$random}};
    R118 = {4{$random}};
    R126 = {1{$random}};
    R131 = {1{$random}};
    R164 = {1{$random}};
    R218 = {1{$random}};
    R228 = {1{$random}};
    R238 = {1{$random}};
    R255 = {2{$random}};
    R261 = {2{$random}};
    R277 = {1{$random}};
    R283 = {1{$random}};
    R289 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T15 | T3;
  assign T3 = T14 ? 1'h1 : T4;
  assign T4 = T13 ? 1'h1 : T5;
  assign T5 = T12 ? 1'h1 : T6;
  assign T6 = T11 ? 1'h1 : T7;
  assign T7 = T10 ? 1'h1 : T8;
  assign T8 = T9 == 3'h3;
  assign T9 = io_in_acquire_bits_union[4'h8:3'h6];
  assign T10 = T9 == 3'h2;
  assign T11 = T9 == 3'h5;
  assign T12 = T9 == 3'h1;
  assign T13 = T9 == 3'h4;
  assign T14 = T9 == 3'h0;
  assign T15 = T18 | T16;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_in_acquire_bits_a_type == 3'h0;
  assign T18 = io_in_acquire_valid ^ 1'h1;
  assign T20 = T21 | reset;
  assign T21 = T70 | T22;
  assign T22 = T23 <= 2'h1;
  assign T23 = T306 + T24;
  assign T24 = {1'h0, T25};
  assign T25 = T26[1'h1:1'h1];
  assign T26 = {T48, T27};
  assign T27 = T28 != 8'h0;
  assign T28 = T29[3'h7:1'h0];
  assign T29 = T46 ? T37 : T30;
  assign T30 = T32 ? T31 : 16'h0;
  assign T31 = io_in_acquire_bits_union[5'h10:1'h1];
  assign T32 = T35 | T33;
  assign T33 = io_in_acquire_bits_is_builtin_type & T34;
  assign T34 = io_in_acquire_bits_a_type == 3'h2;
  assign T35 = io_in_acquire_bits_is_builtin_type & T36;
  assign T36 = io_in_acquire_bits_a_type == 3'h3;
  assign T37 = T38;
  assign T38 = {T44, T39};
  assign T39 = 8'h0 - T302;
  assign T302 = {7'h0, T40};
  assign T40 = T41[1'h0:1'h0];
  assign T41 = 1'h1 << T42;
  assign T42 = T43[2'h3:2'h3];
  assign T43 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T44 = 8'h0 - T303;
  assign T303 = {7'h0, T45};
  assign T45 = T41[1'h1:1'h1];
  assign T46 = io_in_acquire_bits_is_builtin_type & T47;
  assign T47 = io_in_acquire_bits_a_type == 3'h4;
  assign T48 = T49 != 8'h0;
  assign T49 = T50[4'hf:4'h8];
  assign T50 = T67 ? T58 : T51;
  assign T51 = T53 ? T52 : 16'h0;
  assign T52 = io_in_acquire_bits_union[5'h10:1'h1];
  assign T53 = T56 | T54;
  assign T54 = io_in_acquire_bits_is_builtin_type & T55;
  assign T55 = io_in_acquire_bits_a_type == 3'h2;
  assign T56 = io_in_acquire_bits_is_builtin_type & T57;
  assign T57 = io_in_acquire_bits_a_type == 3'h3;
  assign T58 = T59;
  assign T59 = {T65, T60};
  assign T60 = 8'h0 - T304;
  assign T304 = {7'h0, T61};
  assign T61 = T62[1'h0:1'h0];
  assign T62 = 1'h1 << T63;
  assign T63 = T64[2'h3:2'h3];
  assign T64 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T65 = 8'h0 - T305;
  assign T305 = {7'h0, T66};
  assign T66 = T62[1'h1:1'h1];
  assign T67 = io_in_acquire_bits_is_builtin_type & T68;
  assign T68 = io_in_acquire_bits_a_type == 3'h4;
  assign T306 = {1'h0, T69};
  assign T69 = T26[1'h0:1'h0];
  assign T70 = T73 | T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = io_in_acquire_bits_a_type == 3'h2;
  assign T73 = io_in_acquire_valid ^ 1'h1;
  assign T74 = T76 & T75;
  assign T75 = io_out_grant_bits_g_type == 4'h4;
  assign T76 = io_out_grant_ready & io_out_grant_valid;
  assign T77 = T78[2'h3:2'h3];
  assign T78 = {io_in_acquire_bits_addr_block, T79};
  assign T79 = {io_in_acquire_bits_addr_beat, T80};
  assign T80 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T81 = T82 & io_out_acquire_ready;
  assign T82 = T17 & io_in_acquire_valid;
  assign io_out_grant_ready = T83;
  assign T83 = T88 & T84;
  assign T84 = T85 | io_in_grant_ready;
  assign T85 = io_out_grant_bits_is_builtin_type ? T87 : T86;
  assign T86 = 4'h0 == io_out_grant_bits_g_type;
  assign T87 = 4'h5 == io_out_grant_bits_g_type;
  assign T88 = R89 ^ 1'h1;
  assign T307 = reset ? 1'h0 : T90;
  assign T90 = T100 ? 1'h0 : T91;
  assign T91 = T92 ? 1'h1 : R89;
  assign T92 = T97 & T93;
  assign T93 = R94 == 1'h1;
  assign T308 = reset ? 1'h0 : T95;
  assign T95 = T97 ? T96 : R94;
  assign T96 = R94 + 1'h1;
  assign T97 = T99 & T98;
  assign T98 = R89 ^ 1'h1;
  assign T99 = io_out_grant_valid & T85;
  assign T100 = io_in_grant_ready & R89;
  assign io_out_acquire_bits_data = T309;
  assign T309 = T101[6'h3f:1'h0];
  assign T101 = R126 ? T313 : T102;
  assign T102 = T115 ? T312 : T103;
  assign T103 = T72 ? T311 : T104;
  assign T104 = T17 ? T310 : io_in_acquire_bits_data;
  assign T310 = {64'h0, T105};
  assign T105 = 64'h0;
  assign T311 = {64'h0, T106};
  assign T106 = T107;
  assign T107 = T111 | T108;
  assign T108 = T110 ? T109 : 64'h0;
  assign T109 = io_in_acquire_bits_data[7'h7f:7'h40];
  assign T110 = T26[1'h1:1'h1];
  assign T111 = T113 ? T112 : 64'h0;
  assign T112 = io_in_acquire_bits_data[6'h3f:1'h0];
  assign T113 = T26[1'h0:1'h0];
  assign T312 = {64'h0, T114};
  assign T114 = 64'h0;
  assign T115 = io_in_acquire_bits_a_type == 3'h1;
  assign T313 = {64'h0, T116};
  assign T116 = T117;
  assign T117 = R118[6'h3f:1'h0];
  assign T119 = T125 ? T314 : T120;
  assign T120 = T121 ? io_in_acquire_bits_data : R118;
  assign T121 = T123 & T122;
  assign T122 = io_in_acquire_bits_a_type == 3'h3;
  assign T123 = io_in_acquire_ready & io_in_acquire_valid;
  assign T314 = {64'h0, T124};
  assign T124 = R118 >> 7'h40;
  assign T125 = R126 & io_out_acquire_ready;
  assign T315 = reset ? 1'h0 : T127;
  assign T127 = T129 ? 1'h0 : T128;
  assign T128 = T121 ? 1'h1 : R126;
  assign T129 = T125 & T130;
  assign T130 = R131 == 1'h1;
  assign T316 = reset ? 1'h0 : T132;
  assign T132 = T125 ? T133 : R131;
  assign T133 = R131 + 1'h1;
  assign io_out_acquire_bits_union = T317;
  assign T317 = T134[4'hb:1'h0];
  assign T134 = R126 ? T323 : T135;
  assign T135 = T115 ? T321 : T136;
  assign T136 = T72 ? T319 : T137;
  assign T137 = T17 ? T318 : io_in_acquire_bits_union;
  assign T318 = {5'h0, T138};
  assign T138 = T139;
  assign T139 = {T142, T140};
  assign T140 = {5'h0, T141};
  assign T141 = io_in_acquire_bits_union[1'h0:1'h0];
  assign T142 = {T144, T143};
  assign T143 = io_in_acquire_bits_union[4'h8:3'h6];
  assign T144 = T145[2'h2:1'h0];
  assign T145 = {io_in_acquire_bits_addr_block, T146};
  assign T146 = {io_in_acquire_bits_addr_beat, T147};
  assign T147 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T319 = {5'h0, T148};
  assign T148 = T320;
  assign T320 = {3'h0, T149};
  assign T149 = {T150, 1'h1};
  assign T150 = T153 | T151;
  assign T151 = T152 ? T49 : 8'h0;
  assign T152 = T26[1'h1:1'h1];
  assign T153 = T154 ? T28 : 8'h0;
  assign T154 = T26[1'h0:1'h0];
  assign T321 = {5'h0, T155};
  assign T155 = T322;
  assign T322 = {3'h0, T156};
  assign T156 = {3'h7, T157};
  assign T157 = {5'h0, T158};
  assign T158 = io_in_acquire_bits_union[1'h0:1'h0];
  assign T323 = {5'h0, T159};
  assign T159 = T324;
  assign T324 = {3'h0, T160};
  assign T160 = {T163, T161};
  assign T161 = T163 != T162;
  assign T162 = 8'hff;
  assign T163 = R164[3'h7:1'h0];
  assign T165 = T125 ? T327 : T166;
  assign T166 = T121 ? T167 : R164;
  assign T167 = T184 ? T175 : T168;
  assign T168 = T170 ? T169 : 16'h0;
  assign T169 = io_in_acquire_bits_union[5'h10:1'h1];
  assign T170 = T173 | T171;
  assign T171 = io_in_acquire_bits_is_builtin_type & T172;
  assign T172 = io_in_acquire_bits_a_type == 3'h2;
  assign T173 = io_in_acquire_bits_is_builtin_type & T174;
  assign T174 = io_in_acquire_bits_a_type == 3'h3;
  assign T175 = T176;
  assign T176 = {T182, T177};
  assign T177 = 8'h0 - T325;
  assign T325 = {7'h0, T178};
  assign T178 = T179[1'h0:1'h0];
  assign T179 = 1'h1 << T180;
  assign T180 = T181[2'h3:2'h3];
  assign T181 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T182 = 8'h0 - T326;
  assign T326 = {7'h0, T183};
  assign T183 = T179[1'h1:1'h1];
  assign T184 = io_in_acquire_bits_is_builtin_type & T185;
  assign T185 = io_in_acquire_bits_a_type == 3'h4;
  assign T327 = {8'h0, T186};
  assign T186 = R164 >> 4'h8;
  assign io_out_acquire_bits_a_type = T187;
  assign T187 = R126 ? T194 : T188;
  assign T188 = T115 ? T193 : T189;
  assign T189 = T72 ? T192 : T190;
  assign T190 = T17 ? T191 : io_in_acquire_bits_a_type;
  assign T191 = 3'h0;
  assign T192 = 3'h2;
  assign T193 = 3'h1;
  assign T194 = 3'h3;
  assign io_out_acquire_bits_is_builtin_type = T195;
  assign T195 = R126 ? T202 : T196;
  assign T196 = T115 ? T201 : T197;
  assign T197 = T72 ? T200 : T198;
  assign T198 = T17 ? T199 : io_in_acquire_bits_is_builtin_type;
  assign T199 = 1'h1;
  assign T200 = 1'h1;
  assign T201 = 1'h1;
  assign T202 = 1'h1;
  assign io_out_acquire_bits_addr_beat = T203;
  assign T203 = R126 ? T216 : T204;
  assign T204 = T115 ? T215 : T205;
  assign T205 = T72 ? T212 : T206;
  assign T206 = T17 ? T207 : T328;
  assign T328 = {1'h0, io_in_acquire_bits_addr_beat};
  assign T207 = T208;
  assign T208 = T209[3'h5:2'h3];
  assign T209 = {io_in_acquire_bits_addr_block, T210};
  assign T210 = {io_in_acquire_bits_addr_beat, T211};
  assign T211 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T212 = T213;
  assign T213 = {io_in_acquire_bits_addr_beat, T329};
  assign T329 = T330 == 1'h0;
  assign T330 = T26[1'h0:1'h0];
  assign T215 = 3'h0;
  assign T216 = T217;
  assign T217 = {R218, R131};
  assign T219 = T121 ? io_in_acquire_bits_addr_beat : R218;
  assign io_out_acquire_bits_client_xact_id = T220;
  assign T220 = R126 ? T227 : T221;
  assign T221 = T115 ? T226 : T222;
  assign T222 = T72 ? T225 : T223;
  assign T223 = T17 ? T224 : io_in_acquire_bits_client_xact_id;
  assign T224 = io_in_acquire_bits_client_xact_id;
  assign T225 = io_in_acquire_bits_client_xact_id;
  assign T226 = io_in_acquire_bits_client_xact_id;
  assign T227 = R228;
  assign T229 = T121 ? io_in_acquire_bits_client_xact_id : R228;
  assign io_out_acquire_bits_addr_block = T230;
  assign T230 = R126 ? T237 : T231;
  assign T231 = T115 ? T236 : T232;
  assign T232 = T72 ? T235 : T233;
  assign T233 = T17 ? T234 : io_in_acquire_bits_addr_block;
  assign T234 = io_in_acquire_bits_addr_block;
  assign T235 = io_in_acquire_bits_addr_block;
  assign T236 = io_in_acquire_bits_addr_block;
  assign T237 = R238;
  assign T239 = T121 ? io_in_acquire_bits_addr_block : R238;
  assign io_out_acquire_valid = T240;
  assign T240 = T242 | T241;
  assign T241 = T82 & ReorderQueue_io_enq_ready;
  assign T242 = R126 | T243;
  assign T243 = T245 & T244;
  assign T244 = T17 ^ 1'h1;
  assign T245 = io_in_acquire_valid & T246;
  assign T246 = T122 ^ 1'h1;
  assign io_in_grant_bits_data = T247;
  assign T247 = R89 ? T252 : T248;
  assign T248 = T75 ? T249 : T331;
  assign T331 = {64'h0, io_out_grant_bits_data};
  assign T249 = T332;
  assign T332 = T250[7'h7f:1'h0];
  assign T250 = io_out_grant_bits_data << T251;
  assign T251 = {ReorderQueue_io_deq_data, 6'h0};
  assign T252 = T253;
  assign T253 = T254;
  assign T254 = {R261, R255};
  assign T256 = T257 ? io_out_grant_bits_data : R255;
  assign T257 = T97 & T258;
  assign T258 = T259[1'h0:1'h0];
  assign T259 = 1'h1 << T260;
  assign T260 = R94;
  assign T262 = T263 ? io_out_grant_bits_data : R261;
  assign T263 = T97 & T264;
  assign T264 = T259[1'h1:1'h1];
  assign io_in_grant_bits_g_type = T265;
  assign T265 = R89 ? T268 : T266;
  assign T266 = T75 ? T267 : io_out_grant_bits_g_type;
  assign T267 = 4'h4;
  assign T268 = 4'h5;
  assign io_in_grant_bits_is_builtin_type = T269;
  assign T269 = R89 ? T272 : T270;
  assign T270 = T75 ? T271 : io_out_grant_bits_is_builtin_type;
  assign T271 = 1'h1;
  assign T272 = 1'h1;
  assign io_in_grant_bits_manager_xact_id = T273;
  assign T273 = R89 ? T276 : T274;
  assign T274 = T75 ? T275 : io_out_grant_bits_manager_xact_id;
  assign T275 = io_out_grant_bits_manager_xact_id;
  assign T276 = R277;
  assign T278 = T92 ? io_out_grant_bits_manager_xact_id : R277;
  assign io_in_grant_bits_client_xact_id = T279;
  assign T279 = R89 ? T282 : T280;
  assign T280 = T75 ? T281 : io_out_grant_bits_client_xact_id;
  assign T281 = io_out_grant_bits_client_xact_id;
  assign T282 = R283;
  assign T284 = T92 ? io_out_grant_bits_client_xact_id : R283;
  assign io_in_grant_bits_addr_beat = T333;
  assign T333 = T285[1'h1:1'h0];
  assign T285 = R89 ? T336 : T286;
  assign T286 = T75 ? T334 : io_out_grant_bits_addr_beat;
  assign T334 = {1'h0, T287};
  assign T287 = T335;
  assign T335 = io_out_grant_bits_addr_beat[1'h1:1'h0];
  assign T336 = {1'h0, T288};
  assign T288 = R289;
  assign T337 = reset ? 2'h0 : T290;
  assign T290 = T100 ? T291 : R289;
  assign T291 = R289 + 2'h1;
  assign io_in_grant_valid = T292;
  assign T292 = R89 | T293;
  assign T293 = io_out_grant_valid & T294;
  assign T294 = T85 ^ 1'h1;
  assign io_in_acquire_ready = T295;
  assign T295 = T301 & T296;
  assign T296 = T298 | T297;
  assign T297 = ReorderQueue_io_enq_ready & io_out_acquire_ready;
  assign T298 = T122 | T299;
  assign T299 = T300 & io_out_acquire_ready;
  assign T300 = T17 ^ 1'h1;
  assign T301 = R126 ^ 1'h1;
  ReorderQueue_0 ReorderQueue(.clk(clk), .reset(reset),
       .io_enq_ready( ReorderQueue_io_enq_ready ),
       .io_enq_valid( T81 ),
       .io_enq_bits_data( T77 ),
       .io_enq_bits_tag( io_in_acquire_bits_client_xact_id ),
       .io_deq_valid( T74 ),
       .io_deq_tag( io_out_grant_bits_client_xact_id ),
       .io_deq_data( ReorderQueue_io_deq_data )
       //.io_deq_matches(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T19 <= 1'b1;
  if(!T20 && T19 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't perform Put wider than outer width");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't perform Get wider than outer width");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      R89 <= 1'h0;
    end else if(T100) begin
      R89 <= 1'h0;
    end else if(T92) begin
      R89 <= 1'h1;
    end
    if(reset) begin
      R94 <= 1'h0;
    end else if(T97) begin
      R94 <= T96;
    end
    if(T125) begin
      R118 <= T314;
    end else if(T121) begin
      R118 <= io_in_acquire_bits_data;
    end
    if(reset) begin
      R126 <= 1'h0;
    end else if(T129) begin
      R126 <= 1'h0;
    end else if(T121) begin
      R126 <= 1'h1;
    end
    if(reset) begin
      R131 <= 1'h0;
    end else if(T125) begin
      R131 <= T133;
    end
    if(T125) begin
      R164 <= T327;
    end else if(T121) begin
      R164 <= T167;
    end
    if(T121) begin
      R218 <= io_in_acquire_bits_addr_beat;
    end
    if(T121) begin
      R228 <= io_in_acquire_bits_client_xact_id;
    end
    if(T121) begin
      R238 <= io_in_acquire_bits_addr_block;
    end
    if(T257) begin
      R255 <= io_out_grant_bits_data;
    end
    if(T263) begin
      R261 <= io_out_grant_bits_data;
    end
    if(T92) begin
      R277 <= io_out_grant_bits_manager_xact_id;
    end
    if(T92) begin
      R283 <= io_out_grant_bits_client_xact_id;
    end
    if(reset) begin
      R289 <= 2'h0;
    end else if(T100) begin
      R289 <= T291;
    end
  end
endmodule

module ReorderQueue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_data_byteOff,
    input  io_enq_bits_data_subblock,
    input [4:0] io_enq_bits_tag,
    input  io_deq_valid,
    input [4:0] io_deq_tag,
    output[2:0] io_deq_data_byteOff,
    output io_deq_data_subblock,
    output io_deq_matches
);

  wire T0;
  wire roq_matches_8;
  wire T1;
  reg  roq_free_8;
  wire T216;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[15:0] T6;
  wire[3:0] T7;
  wire[3:0] roq_enq_addr;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  reg  roq_free_7;
  wire T217;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[15:0] T21;
  wire[3:0] T22;
  wire[3:0] roq_deq_addr;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  wire roq_matches_7;
  wire T30;
  wire T31;
  reg [4:0] roq_tags_7;
  wire[4:0] T32;
  wire T33;
  wire T34;
  wire[15:0] T35;
  wire[3:0] T36;
  wire roq_matches_6;
  wire T37;
  wire T38;
  reg [4:0] roq_tags_6;
  wire[4:0] T39;
  wire T40;
  wire T41;
  wire roq_matches_5;
  wire T42;
  wire T43;
  reg [4:0] roq_tags_5;
  wire[4:0] T44;
  wire T45;
  wire T46;
  wire roq_matches_4;
  wire T47;
  wire T48;
  reg [4:0] roq_tags_4;
  wire[4:0] T49;
  wire T50;
  wire T51;
  wire roq_matches_3;
  wire T52;
  wire T53;
  reg [4:0] roq_tags_3;
  wire[4:0] T54;
  wire T55;
  wire T56;
  wire roq_matches_2;
  wire T57;
  wire T58;
  reg [4:0] roq_tags_2;
  wire[4:0] T59;
  wire T60;
  wire T61;
  wire roq_matches_1;
  wire T62;
  wire T63;
  reg [4:0] roq_tags_1;
  wire[4:0] T64;
  wire T65;
  wire T66;
  wire roq_matches_0;
  wire T67;
  wire T68;
  reg [4:0] roq_tags_0;
  wire[4:0] T69;
  wire T70;
  wire T71;
  reg  roq_free_6;
  wire T218;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg  roq_free_5;
  wire T219;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  reg  roq_free_4;
  wire T220;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg  roq_free_3;
  wire T221;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  reg  roq_free_2;
  wire T222;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  reg  roq_free_1;
  wire T223;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg  roq_free_0;
  wire T224;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  reg [4:0] roq_tags_8;
  wire[4:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg  roq_data_0_subblock;
  wire T132;
  wire T133;
  wire T134;
  wire[15:0] T135;
  wire[3:0] T136;
  reg  roq_data_1_subblock;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire[3:0] T141;
  wire T142;
  reg  roq_data_2_subblock;
  wire T143;
  wire T144;
  wire T145;
  reg  roq_data_3_subblock;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg  roq_data_4_subblock;
  wire T153;
  wire T154;
  wire T155;
  reg  roq_data_5_subblock;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  reg  roq_data_6_subblock;
  wire T161;
  wire T162;
  wire T163;
  reg  roq_data_7_subblock;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  reg  roq_data_8_subblock;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire[2:0] T174;
  wire[2:0] T175;
  wire[2:0] T176;
  wire[2:0] T177;
  reg [2:0] roq_data_0_byteOff;
  wire[2:0] T178;
  wire T179;
  reg [2:0] roq_data_1_byteOff;
  wire[2:0] T180;
  wire T181;
  wire T182;
  wire[2:0] T183;
  reg [2:0] roq_data_2_byteOff;
  wire[2:0] T184;
  wire T185;
  reg [2:0] roq_data_3_byteOff;
  wire[2:0] T186;
  wire T187;
  wire T188;
  wire T189;
  wire[2:0] T190;
  wire[2:0] T191;
  reg [2:0] roq_data_4_byteOff;
  wire[2:0] T192;
  wire T193;
  reg [2:0] roq_data_5_byteOff;
  wire[2:0] T194;
  wire T195;
  wire T196;
  wire[2:0] T197;
  reg [2:0] roq_data_6_byteOff;
  wire[2:0] T198;
  wire T199;
  reg [2:0] roq_data_7_byteOff;
  wire[2:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  reg [2:0] roq_data_8_byteOff;
  wire[2:0] T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    roq_free_8 = {1{$random}};
    roq_free_7 = {1{$random}};
    roq_tags_7 = {1{$random}};
    roq_tags_6 = {1{$random}};
    roq_tags_5 = {1{$random}};
    roq_tags_4 = {1{$random}};
    roq_tags_3 = {1{$random}};
    roq_tags_2 = {1{$random}};
    roq_tags_1 = {1{$random}};
    roq_tags_0 = {1{$random}};
    roq_free_6 = {1{$random}};
    roq_free_5 = {1{$random}};
    roq_free_4 = {1{$random}};
    roq_free_3 = {1{$random}};
    roq_free_2 = {1{$random}};
    roq_free_1 = {1{$random}};
    roq_free_0 = {1{$random}};
    roq_tags_8 = {1{$random}};
    roq_data_0_subblock = {1{$random}};
    roq_data_1_subblock = {1{$random}};
    roq_data_2_subblock = {1{$random}};
    roq_data_3_subblock = {1{$random}};
    roq_data_4_subblock = {1{$random}};
    roq_data_5_subblock = {1{$random}};
    roq_data_6_subblock = {1{$random}};
    roq_data_7_subblock = {1{$random}};
    roq_data_8_subblock = {1{$random}};
    roq_data_0_byteOff = {1{$random}};
    roq_data_1_byteOff = {1{$random}};
    roq_data_2_byteOff = {1{$random}};
    roq_data_3_byteOff = {1{$random}};
    roq_data_4_byteOff = {1{$random}};
    roq_data_5_byteOff = {1{$random}};
    roq_data_6_byteOff = {1{$random}};
    roq_data_7_byteOff = {1{$random}};
    roq_data_8_byteOff = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_deq_matches = T0;
  assign T0 = T121 | roq_matches_8;
  assign roq_matches_8 = T117 & T1;
  assign T1 = roq_free_8 ^ 1'h1;
  assign T216 = reset ? 1'h1 : T2;
  assign T2 = T115 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : roq_free_8;
  assign T4 = T114 & T5;
  assign T5 = T6[4'h8:4'h8];
  assign T6 = 1'h1 << T7;
  assign T7 = roq_enq_addr;
  assign roq_enq_addr = roq_free_0 ? 4'h0 : T8;
  assign T8 = roq_free_1 ? 4'h1 : T9;
  assign T9 = roq_free_2 ? 4'h2 : T10;
  assign T10 = roq_free_3 ? 4'h3 : T11;
  assign T11 = roq_free_4 ? 4'h4 : T12;
  assign T12 = roq_free_5 ? 4'h5 : T13;
  assign T13 = roq_free_6 ? 4'h6 : T14;
  assign T14 = roq_free_7 ? 4'h7 : 4'h8;
  assign T217 = reset ? 1'h1 : T15;
  assign T15 = T19 ? 1'h1 : T16;
  assign T16 = T17 ? 1'h0 : roq_free_7;
  assign T17 = T114 & T18;
  assign T18 = T6[3'h7:3'h7];
  assign T19 = io_deq_valid & T20;
  assign T20 = T21[3'h7:3'h7];
  assign T21 = 1'h1 << T22;
  assign T22 = roq_deq_addr;
  assign roq_deq_addr = roq_matches_0 ? 4'h0 : T23;
  assign T23 = roq_matches_1 ? 4'h1 : T24;
  assign T24 = roq_matches_2 ? 4'h2 : T25;
  assign T25 = roq_matches_3 ? 4'h3 : T26;
  assign T26 = roq_matches_4 ? 4'h4 : T27;
  assign T27 = roq_matches_5 ? 4'h5 : T28;
  assign T28 = roq_matches_6 ? 4'h6 : T29;
  assign T29 = roq_matches_7 ? 4'h7 : 4'h8;
  assign roq_matches_7 = T31 & T30;
  assign T30 = roq_free_7 ^ 1'h1;
  assign T31 = roq_tags_7 == io_deq_tag;
  assign T32 = T33 ? io_enq_bits_tag : roq_tags_7;
  assign T33 = T114 & T34;
  assign T34 = T35[3'h7:3'h7];
  assign T35 = 1'h1 << T36;
  assign T36 = roq_enq_addr;
  assign roq_matches_6 = T38 & T37;
  assign T37 = roq_free_6 ^ 1'h1;
  assign T38 = roq_tags_6 == io_deq_tag;
  assign T39 = T40 ? io_enq_bits_tag : roq_tags_6;
  assign T40 = T114 & T41;
  assign T41 = T35[3'h6:3'h6];
  assign roq_matches_5 = T43 & T42;
  assign T42 = roq_free_5 ^ 1'h1;
  assign T43 = roq_tags_5 == io_deq_tag;
  assign T44 = T45 ? io_enq_bits_tag : roq_tags_5;
  assign T45 = T114 & T46;
  assign T46 = T35[3'h5:3'h5];
  assign roq_matches_4 = T48 & T47;
  assign T47 = roq_free_4 ^ 1'h1;
  assign T48 = roq_tags_4 == io_deq_tag;
  assign T49 = T50 ? io_enq_bits_tag : roq_tags_4;
  assign T50 = T114 & T51;
  assign T51 = T35[3'h4:3'h4];
  assign roq_matches_3 = T53 & T52;
  assign T52 = roq_free_3 ^ 1'h1;
  assign T53 = roq_tags_3 == io_deq_tag;
  assign T54 = T55 ? io_enq_bits_tag : roq_tags_3;
  assign T55 = T114 & T56;
  assign T56 = T35[2'h3:2'h3];
  assign roq_matches_2 = T58 & T57;
  assign T57 = roq_free_2 ^ 1'h1;
  assign T58 = roq_tags_2 == io_deq_tag;
  assign T59 = T60 ? io_enq_bits_tag : roq_tags_2;
  assign T60 = T114 & T61;
  assign T61 = T35[2'h2:2'h2];
  assign roq_matches_1 = T63 & T62;
  assign T62 = roq_free_1 ^ 1'h1;
  assign T63 = roq_tags_1 == io_deq_tag;
  assign T64 = T65 ? io_enq_bits_tag : roq_tags_1;
  assign T65 = T114 & T66;
  assign T66 = T35[1'h1:1'h1];
  assign roq_matches_0 = T68 & T67;
  assign T67 = roq_free_0 ^ 1'h1;
  assign T68 = roq_tags_0 == io_deq_tag;
  assign T69 = T70 ? io_enq_bits_tag : roq_tags_0;
  assign T70 = T114 & T71;
  assign T71 = T35[1'h0:1'h0];
  assign T218 = reset ? 1'h1 : T72;
  assign T72 = T76 ? 1'h1 : T73;
  assign T73 = T74 ? 1'h0 : roq_free_6;
  assign T74 = T114 & T75;
  assign T75 = T6[3'h6:3'h6];
  assign T76 = io_deq_valid & T77;
  assign T77 = T21[3'h6:3'h6];
  assign T219 = reset ? 1'h1 : T78;
  assign T78 = T82 ? 1'h1 : T79;
  assign T79 = T80 ? 1'h0 : roq_free_5;
  assign T80 = T114 & T81;
  assign T81 = T6[3'h5:3'h5];
  assign T82 = io_deq_valid & T83;
  assign T83 = T21[3'h5:3'h5];
  assign T220 = reset ? 1'h1 : T84;
  assign T84 = T88 ? 1'h1 : T85;
  assign T85 = T86 ? 1'h0 : roq_free_4;
  assign T86 = T114 & T87;
  assign T87 = T6[3'h4:3'h4];
  assign T88 = io_deq_valid & T89;
  assign T89 = T21[3'h4:3'h4];
  assign T221 = reset ? 1'h1 : T90;
  assign T90 = T94 ? 1'h1 : T91;
  assign T91 = T92 ? 1'h0 : roq_free_3;
  assign T92 = T114 & T93;
  assign T93 = T6[2'h3:2'h3];
  assign T94 = io_deq_valid & T95;
  assign T95 = T21[2'h3:2'h3];
  assign T222 = reset ? 1'h1 : T96;
  assign T96 = T100 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : roq_free_2;
  assign T98 = T114 & T99;
  assign T99 = T6[2'h2:2'h2];
  assign T100 = io_deq_valid & T101;
  assign T101 = T21[2'h2:2'h2];
  assign T223 = reset ? 1'h1 : T102;
  assign T102 = T106 ? 1'h1 : T103;
  assign T103 = T104 ? 1'h0 : roq_free_1;
  assign T104 = T114 & T105;
  assign T105 = T6[1'h1:1'h1];
  assign T106 = io_deq_valid & T107;
  assign T107 = T21[1'h1:1'h1];
  assign T224 = reset ? 1'h1 : T108;
  assign T108 = T112 ? 1'h1 : T109;
  assign T109 = T110 ? 1'h0 : roq_free_0;
  assign T110 = T114 & T111;
  assign T111 = T6[1'h0:1'h0];
  assign T112 = io_deq_valid & T113;
  assign T113 = T21[1'h0:1'h0];
  assign T114 = io_enq_valid & io_enq_ready;
  assign T115 = io_deq_valid & T116;
  assign T116 = T21[4'h8:4'h8];
  assign T117 = roq_tags_8 == io_deq_tag;
  assign T118 = T119 ? io_enq_bits_tag : roq_tags_8;
  assign T119 = T114 & T120;
  assign T120 = T35[4'h8:4'h8];
  assign T121 = T122 | roq_matches_7;
  assign T122 = T123 | roq_matches_6;
  assign T123 = T124 | roq_matches_5;
  assign T124 = T125 | roq_matches_4;
  assign T125 = T126 | roq_matches_3;
  assign T126 = T127 | roq_matches_2;
  assign T127 = roq_matches_0 | roq_matches_1;
  assign io_deq_data_subblock = T128;
  assign T128 = T173 ? roq_data_8_subblock : T129;
  assign T129 = T169 ? T151 : T130;
  assign T130 = T150 ? T142 : T131;
  assign T131 = T140 ? roq_data_1_subblock : roq_data_0_subblock;
  assign T132 = T133 ? io_enq_bits_data_subblock : roq_data_0_subblock;
  assign T133 = T114 & T134;
  assign T134 = T135[1'h0:1'h0];
  assign T135 = 1'h1 << T136;
  assign T136 = roq_enq_addr;
  assign T137 = T138 ? io_enq_bits_data_subblock : roq_data_1_subblock;
  assign T138 = T114 & T139;
  assign T139 = T135[1'h1:1'h1];
  assign T140 = T141[1'h0:1'h0];
  assign T141 = roq_deq_addr;
  assign T142 = T149 ? roq_data_3_subblock : roq_data_2_subblock;
  assign T143 = T144 ? io_enq_bits_data_subblock : roq_data_2_subblock;
  assign T144 = T114 & T145;
  assign T145 = T135[2'h2:2'h2];
  assign T146 = T147 ? io_enq_bits_data_subblock : roq_data_3_subblock;
  assign T147 = T114 & T148;
  assign T148 = T135[2'h3:2'h3];
  assign T149 = T141[1'h0:1'h0];
  assign T150 = T141[1'h1:1'h1];
  assign T151 = T168 ? T160 : T152;
  assign T152 = T159 ? roq_data_5_subblock : roq_data_4_subblock;
  assign T153 = T154 ? io_enq_bits_data_subblock : roq_data_4_subblock;
  assign T154 = T114 & T155;
  assign T155 = T135[3'h4:3'h4];
  assign T156 = T157 ? io_enq_bits_data_subblock : roq_data_5_subblock;
  assign T157 = T114 & T158;
  assign T158 = T135[3'h5:3'h5];
  assign T159 = T141[1'h0:1'h0];
  assign T160 = T167 ? roq_data_7_subblock : roq_data_6_subblock;
  assign T161 = T162 ? io_enq_bits_data_subblock : roq_data_6_subblock;
  assign T162 = T114 & T163;
  assign T163 = T135[3'h6:3'h6];
  assign T164 = T165 ? io_enq_bits_data_subblock : roq_data_7_subblock;
  assign T165 = T114 & T166;
  assign T166 = T135[3'h7:3'h7];
  assign T167 = T141[1'h0:1'h0];
  assign T168 = T141[1'h1:1'h1];
  assign T169 = T141[2'h2:2'h2];
  assign T170 = T171 ? io_enq_bits_data_subblock : roq_data_8_subblock;
  assign T171 = T114 & T172;
  assign T172 = T135[4'h8:4'h8];
  assign T173 = T141[2'h3:2'h3];
  assign io_deq_data_byteOff = T174;
  assign T174 = T207 ? roq_data_8_byteOff : T175;
  assign T175 = T204 ? T190 : T176;
  assign T176 = T189 ? T183 : T177;
  assign T177 = T182 ? roq_data_1_byteOff : roq_data_0_byteOff;
  assign T178 = T179 ? io_enq_bits_data_byteOff : roq_data_0_byteOff;
  assign T179 = T114 & T134;
  assign T180 = T181 ? io_enq_bits_data_byteOff : roq_data_1_byteOff;
  assign T181 = T114 & T139;
  assign T182 = T141[1'h0:1'h0];
  assign T183 = T188 ? roq_data_3_byteOff : roq_data_2_byteOff;
  assign T184 = T185 ? io_enq_bits_data_byteOff : roq_data_2_byteOff;
  assign T185 = T114 & T145;
  assign T186 = T187 ? io_enq_bits_data_byteOff : roq_data_3_byteOff;
  assign T187 = T114 & T148;
  assign T188 = T141[1'h0:1'h0];
  assign T189 = T141[1'h1:1'h1];
  assign T190 = T203 ? T197 : T191;
  assign T191 = T196 ? roq_data_5_byteOff : roq_data_4_byteOff;
  assign T192 = T193 ? io_enq_bits_data_byteOff : roq_data_4_byteOff;
  assign T193 = T114 & T155;
  assign T194 = T195 ? io_enq_bits_data_byteOff : roq_data_5_byteOff;
  assign T195 = T114 & T158;
  assign T196 = T141[1'h0:1'h0];
  assign T197 = T202 ? roq_data_7_byteOff : roq_data_6_byteOff;
  assign T198 = T199 ? io_enq_bits_data_byteOff : roq_data_6_byteOff;
  assign T199 = T114 & T163;
  assign T200 = T201 ? io_enq_bits_data_byteOff : roq_data_7_byteOff;
  assign T201 = T114 & T166;
  assign T202 = T141[1'h0:1'h0];
  assign T203 = T141[1'h1:1'h1];
  assign T204 = T141[2'h2:2'h2];
  assign T205 = T206 ? io_enq_bits_data_byteOff : roq_data_8_byteOff;
  assign T206 = T114 & T172;
  assign T207 = T141[2'h3:2'h3];
  assign io_enq_ready = T208;
  assign T208 = T209 | roq_free_8;
  assign T209 = T210 | roq_free_7;
  assign T210 = T211 | roq_free_6;
  assign T211 = T212 | roq_free_5;
  assign T212 = T213 | roq_free_4;
  assign T213 = T214 | roq_free_3;
  assign T214 = T215 | roq_free_2;
  assign T215 = roq_free_0 | roq_free_1;

  always @(posedge clk) begin
    if(reset) begin
      roq_free_8 <= 1'h1;
    end else if(T115) begin
      roq_free_8 <= 1'h1;
    end else if(T4) begin
      roq_free_8 <= 1'h0;
    end
    if(reset) begin
      roq_free_7 <= 1'h1;
    end else if(T19) begin
      roq_free_7 <= 1'h1;
    end else if(T17) begin
      roq_free_7 <= 1'h0;
    end
    if(T33) begin
      roq_tags_7 <= io_enq_bits_tag;
    end
    if(T40) begin
      roq_tags_6 <= io_enq_bits_tag;
    end
    if(T45) begin
      roq_tags_5 <= io_enq_bits_tag;
    end
    if(T50) begin
      roq_tags_4 <= io_enq_bits_tag;
    end
    if(T55) begin
      roq_tags_3 <= io_enq_bits_tag;
    end
    if(T60) begin
      roq_tags_2 <= io_enq_bits_tag;
    end
    if(T65) begin
      roq_tags_1 <= io_enq_bits_tag;
    end
    if(T70) begin
      roq_tags_0 <= io_enq_bits_tag;
    end
    if(reset) begin
      roq_free_6 <= 1'h1;
    end else if(T76) begin
      roq_free_6 <= 1'h1;
    end else if(T74) begin
      roq_free_6 <= 1'h0;
    end
    if(reset) begin
      roq_free_5 <= 1'h1;
    end else if(T82) begin
      roq_free_5 <= 1'h1;
    end else if(T80) begin
      roq_free_5 <= 1'h0;
    end
    if(reset) begin
      roq_free_4 <= 1'h1;
    end else if(T88) begin
      roq_free_4 <= 1'h1;
    end else if(T86) begin
      roq_free_4 <= 1'h0;
    end
    if(reset) begin
      roq_free_3 <= 1'h1;
    end else if(T94) begin
      roq_free_3 <= 1'h1;
    end else if(T92) begin
      roq_free_3 <= 1'h0;
    end
    if(reset) begin
      roq_free_2 <= 1'h1;
    end else if(T100) begin
      roq_free_2 <= 1'h1;
    end else if(T98) begin
      roq_free_2 <= 1'h0;
    end
    if(reset) begin
      roq_free_1 <= 1'h1;
    end else if(T106) begin
      roq_free_1 <= 1'h1;
    end else if(T104) begin
      roq_free_1 <= 1'h0;
    end
    if(reset) begin
      roq_free_0 <= 1'h1;
    end else if(T112) begin
      roq_free_0 <= 1'h1;
    end else if(T110) begin
      roq_free_0 <= 1'h0;
    end
    if(T119) begin
      roq_tags_8 <= io_enq_bits_tag;
    end
    if(T133) begin
      roq_data_0_subblock <= io_enq_bits_data_subblock;
    end
    if(T138) begin
      roq_data_1_subblock <= io_enq_bits_data_subblock;
    end
    if(T144) begin
      roq_data_2_subblock <= io_enq_bits_data_subblock;
    end
    if(T147) begin
      roq_data_3_subblock <= io_enq_bits_data_subblock;
    end
    if(T154) begin
      roq_data_4_subblock <= io_enq_bits_data_subblock;
    end
    if(T157) begin
      roq_data_5_subblock <= io_enq_bits_data_subblock;
    end
    if(T162) begin
      roq_data_6_subblock <= io_enq_bits_data_subblock;
    end
    if(T165) begin
      roq_data_7_subblock <= io_enq_bits_data_subblock;
    end
    if(T171) begin
      roq_data_8_subblock <= io_enq_bits_data_subblock;
    end
    if(T179) begin
      roq_data_0_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T181) begin
      roq_data_1_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T185) begin
      roq_data_2_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T187) begin
      roq_data_3_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T193) begin
      roq_data_4_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T195) begin
      roq_data_5_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T199) begin
      roq_data_6_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T201) begin
      roq_data_7_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T206) begin
      roq_data_8_byteOff <= io_enq_bits_data_byteOff;
    end
  end
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_addr_beat,
    input [3:0] io_in_1_bits_client_xact_id,
    input  io_in_1_bits_manager_xact_id,
    input  io_in_1_bits_is_builtin_type,
    input [3:0] io_in_1_bits_g_type,
    input [63:0] io_in_1_bits_data,
    input  io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_addr_beat,
    input [3:0] io_in_0_bits_client_xact_id,
    input  io_in_0_bits_manager_xact_id,
    input  io_in_0_bits_is_builtin_type,
    input [3:0] io_in_0_bits_g_type,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[2:0] io_out_bits_addr_beat,
    output[3:0] io_out_bits_client_xact_id,
    output io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[63:0] io_out_bits_data,
    output io_out_bits_client_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire[63:0] T2;
  wire[3:0] T3;
  wire T4;
  wire T5;
  wire[3:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_client_id = T0;
  assign T0 = T1 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T1 = chosen;
  assign io_out_bits_data = T2;
  assign T2 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_g_type = T3;
  assign T3 = T1 ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign io_out_bits_is_builtin_type = T4;
  assign T4 = T1 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign io_out_bits_manager_xact_id = T5;
  assign T5 = T1 ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign io_out_bits_client_xact_id = T6;
  assign T6 = T1 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_beat = T7;
  assign T7 = T1 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module NastiIOTileLinkIOConverter(input clk, input reset,
    output io_tl_acquire_ready,
    input  io_tl_acquire_valid,
    input [25:0] io_tl_acquire_bits_addr_block,
    input [3:0] io_tl_acquire_bits_client_xact_id,
    input [2:0] io_tl_acquire_bits_addr_beat,
    input  io_tl_acquire_bits_is_builtin_type,
    input [2:0] io_tl_acquire_bits_a_type,
    input [11:0] io_tl_acquire_bits_union,
    input [63:0] io_tl_acquire_bits_data,
    input  io_tl_grant_ready,
    output io_tl_grant_valid,
    output[2:0] io_tl_grant_bits_addr_beat,
    output[3:0] io_tl_grant_bits_client_xact_id,
    output io_tl_grant_bits_manager_xact_id,
    output io_tl_grant_bits_is_builtin_type,
    output[3:0] io_tl_grant_bits_g_type,
    output[63:0] io_tl_grant_bits_data,
    input  io_nasti_aw_ready,
    output io_nasti_aw_valid,
    output[31:0] io_nasti_aw_bits_addr,
    output[7:0] io_nasti_aw_bits_len,
    output[2:0] io_nasti_aw_bits_size,
    output[1:0] io_nasti_aw_bits_burst,
    output io_nasti_aw_bits_lock,
    output[3:0] io_nasti_aw_bits_cache,
    output[2:0] io_nasti_aw_bits_prot,
    output[3:0] io_nasti_aw_bits_qos,
    output[3:0] io_nasti_aw_bits_region,
    output[4:0] io_nasti_aw_bits_id,
    output io_nasti_aw_bits_user,
    input  io_nasti_w_ready,
    output io_nasti_w_valid,
    output[63:0] io_nasti_w_bits_data,
    output io_nasti_w_bits_last,
    output[7:0] io_nasti_w_bits_strb,
    output io_nasti_w_bits_user,
    output io_nasti_b_ready,
    input  io_nasti_b_valid,
    input [1:0] io_nasti_b_bits_resp,
    input [4:0] io_nasti_b_bits_id,
    input  io_nasti_b_bits_user,
    input  io_nasti_ar_ready,
    output io_nasti_ar_valid,
    output[31:0] io_nasti_ar_bits_addr,
    output[7:0] io_nasti_ar_bits_len,
    output[2:0] io_nasti_ar_bits_size,
    output[1:0] io_nasti_ar_bits_burst,
    output io_nasti_ar_bits_lock,
    output[3:0] io_nasti_ar_bits_cache,
    output[2:0] io_nasti_ar_bits_prot,
    output[3:0] io_nasti_ar_bits_qos,
    output[3:0] io_nasti_ar_bits_region,
    output[4:0] io_nasti_ar_bits_id,
    output io_nasti_ar_bits_user,
    output io_nasti_r_ready,
    input  io_nasti_r_valid,
    input [1:0] io_nasti_r_bits_resp,
    input [63:0] io_nasti_r_bits_data,
    input  io_nasti_r_bits_last,
    input [4:0] io_nasti_r_bits_id,
    input  io_nasti_r_bits_user
);

  wire[63:0] T0;
  wire[63:0] T134;
  wire[126:0] r_aligned_data;
  wire[126:0] T135;
  wire[126:0] T1;
  wire[5:0] T2;
  wire[3:0] T3;
  wire[3:0] T136;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[3:0] T7;
  wire[3:0] T137;
  wire[2:0] T8;
  reg [2:0] tl_cnt_in;
  wire[2:0] T138;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[63:0] T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  wire[3:0] T20;
  wire[3:0] T139;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire nasti_wrap_out;
  wire T24;
  reg [2:0] nasti_cnt_out;
  wire[2:0] T140;
  wire[2:0] T25;
  wire[2:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire is_subblock;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[2:0] T36;
  wire T37;
  wire get_valid;
  wire T38;
  wire has_data;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[4:0] T45;
  wire[4:0] T141;
  wire[3:0] T46;
  wire[3:0] T47;
  wire[2:0] T48;
  wire[3:0] T49;
  wire T50;
  wire[1:0] T51;
  wire[2:0] T52;
  wire[2:0] T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire[2:0] T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire[2:0] T60;
  wire T61;
  wire[2:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire[7:0] T69;
  wire[7:0] T142;
  wire[2:0] T70;
  wire[31:0] T71;
  wire[31:0] T72;
  wire[5:0] T73;
  wire[2:0] T74;
  wire T75;
  wire T76;
  wire[7:0] T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T143;
  wire T88;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire tl_wrap_out;
  wire T98;
  reg [2:0] tl_cnt_out;
  wire[2:0] T144;
  wire[2:0] T99;
  wire[2:0] T100;
  wire T101;
  wire is_multibeat;
  wire T102;
  wire T103;
  wire[63:0] T104;
  wire T105;
  wire aw_ready;
  reg  w_inflight;
  wire T145;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire put_valid;
  wire T113;
  wire[4:0] T114;
  wire[4:0] T146;
  wire[3:0] T115;
  wire[3:0] T116;
  wire[2:0] T117;
  wire[3:0] T118;
  wire T119;
  wire[1:0] T120;
  wire[2:0] T121;
  wire[7:0] T122;
  wire[7:0] T147;
  wire[2:0] T123;
  wire[31:0] T124;
  wire[31:0] T125;
  wire[5:0] T126;
  wire[2:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire roq_io_enq_ready;
  wire[2:0] roq_io_deq_data_byteOff;
  wire roq_io_deq_data_subblock;
  wire gnt_arb_io_in_1_ready;
  wire gnt_arb_io_in_0_ready;
  wire gnt_arb_io_out_valid;
  wire[2:0] gnt_arb_io_out_bits_addr_beat;
  wire[3:0] gnt_arb_io_out_bits_client_xact_id;
  wire gnt_arb_io_out_bits_manager_xact_id;
  wire gnt_arb_io_out_bits_is_builtin_type;
  wire[3:0] gnt_arb_io_out_bits_g_type;
  wire[63:0] gnt_arb_io_out_bits_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    tl_cnt_in = {1{$random}};
    nasti_cnt_out = {1{$random}};
    tl_cnt_out = {1{$random}};
    w_inflight = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T134;
  assign T134 = r_aligned_data[6'h3f:1'h0];
  assign r_aligned_data = roq_io_deq_data_subblock ? T1 : T135;
  assign T135 = {63'h0, io_nasti_r_bits_data};
  assign T1 = io_nasti_r_bits_data << T2;
  assign T2 = {roq_io_deq_data_byteOff, 3'h0};
  assign T3 = T136;
  assign T136 = {1'h0, T4};
  assign T4 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T5 = 1'h1;
  assign T6 = 1'h0;
  assign T7 = T137;
  assign T137 = io_nasti_r_bits_id[2'h3:1'h0];
  assign T8 = tl_cnt_in;
  assign T138 = reset ? 3'h0 : T9;
  assign T9 = T11 ? T10 : tl_cnt_in;
  assign T10 = tl_cnt_in + 3'h1;
  assign T11 = T15 & T12;
  assign T12 = io_tl_grant_bits_is_builtin_type ? T14 : T13;
  assign T13 = 4'h0 == io_tl_grant_bits_g_type;
  assign T14 = 4'h5 == io_tl_grant_bits_g_type;
  assign T15 = io_tl_grant_ready & io_tl_grant_valid;
  assign T16 = 64'h0;
  assign T17 = 4'h3;
  assign T18 = 1'h1;
  assign T19 = 1'h0;
  assign T20 = T139;
  assign T139 = io_nasti_b_bits_id[2'h3:1'h0];
  assign T21 = 3'h0;
  assign T22 = T30 & T23;
  assign T23 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign nasti_wrap_out = T27 & T24;
  assign T24 = nasti_cnt_out == 3'h7;
  assign T140 = reset ? 3'h0 : T25;
  assign T25 = T27 ? T26 : nasti_cnt_out;
  assign T26 = nasti_cnt_out + 3'h1;
  assign T27 = T29 & T28;
  assign T28 = roq_io_deq_data_subblock ^ 1'h1;
  assign T29 = io_nasti_r_ready & io_nasti_r_valid;
  assign T30 = io_nasti_r_ready & io_nasti_r_valid;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T31;
  assign T31 = T33 | T32;
  assign T32 = 3'h4 == io_tl_acquire_bits_a_type;
  assign T33 = T35 | T34;
  assign T34 = 3'h0 == io_tl_acquire_bits_a_type;
  assign T35 = 3'h2 == io_tl_acquire_bits_a_type;
  assign T36 = io_tl_acquire_bits_union[4'hb:4'h9];
  assign T37 = get_valid & io_nasti_ar_ready;
  assign get_valid = io_tl_acquire_valid & T38;
  assign T38 = has_data ^ 1'h1;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T39;
  assign T39 = T41 | T40;
  assign T40 = 3'h4 == io_tl_acquire_bits_a_type;
  assign T41 = T43 | T42;
  assign T42 = 3'h3 == io_tl_acquire_bits_a_type;
  assign T43 = 3'h2 == io_tl_acquire_bits_a_type;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign io_nasti_ar_bits_user = T44;
  assign T44 = 1'h0;
  assign io_nasti_ar_bits_id = T45;
  assign T45 = T141;
  assign T141 = {1'h0, io_tl_acquire_bits_client_xact_id};
  assign io_nasti_ar_bits_region = T46;
  assign T46 = 4'h0;
  assign io_nasti_ar_bits_qos = T47;
  assign T47 = 4'h0;
  assign io_nasti_ar_bits_prot = T48;
  assign T48 = 3'h0;
  assign io_nasti_ar_bits_cache = T49;
  assign T49 = 4'h0;
  assign io_nasti_ar_bits_lock = T50;
  assign T50 = 1'h0;
  assign io_nasti_ar_bits_burst = T51;
  assign T51 = 2'h1;
  assign io_nasti_ar_bits_size = T52;
  assign T52 = T53;
  assign T53 = is_subblock ? T54 : 3'h3;
  assign T54 = T68 ? 3'h0 : T55;
  assign T55 = T67 ? 3'h0 : T56;
  assign T56 = T66 ? 3'h1 : T57;
  assign T57 = T65 ? 3'h1 : T58;
  assign T58 = T64 ? 3'h2 : T59;
  assign T59 = T63 ? 3'h3 : T60;
  assign T60 = T61 ? 3'h3 : 3'h7;
  assign T61 = T62 == 3'h7;
  assign T62 = io_tl_acquire_bits_union[4'h8:3'h6];
  assign T63 = T62 == 3'h3;
  assign T64 = T62 == 3'h2;
  assign T65 = T62 == 3'h5;
  assign T66 = T62 == 3'h1;
  assign T67 = T62 == 3'h4;
  assign T68 = T62 == 3'h0;
  assign io_nasti_ar_bits_len = T69;
  assign T69 = T142;
  assign T142 = {5'h0, T70};
  assign T70 = is_subblock ? 3'h0 : 3'h7;
  assign io_nasti_ar_bits_addr = T71;
  assign T71 = T72;
  assign T72 = {io_tl_acquire_bits_addr_block, T73};
  assign T73 = {io_tl_acquire_bits_addr_beat, T74};
  assign T74 = io_tl_acquire_bits_union[4'hb:4'h9];
  assign io_nasti_ar_valid = T75;
  assign T75 = get_valid & roq_io_enq_ready;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_w_bits_user = T76;
  assign T76 = 1'h0;
  assign io_nasti_w_bits_strb = T77;
  assign T77 = T78;
  assign T78 = T92 ? T86 : T79;
  assign T79 = T81 ? T80 : 8'h0;
  assign T80 = io_tl_acquire_bits_union[4'h8:1'h1];
  assign T81 = T84 | T82;
  assign T82 = io_tl_acquire_bits_is_builtin_type & T83;
  assign T83 = io_tl_acquire_bits_a_type == 3'h2;
  assign T84 = io_tl_acquire_bits_is_builtin_type & T85;
  assign T85 = io_tl_acquire_bits_a_type == 3'h3;
  assign T86 = T87;
  assign T87 = 8'h0 - T143;
  assign T143 = {7'h0, T88};
  assign T88 = 1'h1;
  assign T92 = io_tl_acquire_bits_is_builtin_type & T93;
  assign T93 = io_tl_acquire_bits_a_type == 3'h4;
  assign io_nasti_w_bits_last = T94;
  assign T94 = T95;
  assign T95 = tl_wrap_out | T96;
  assign T96 = T97 & is_subblock;
  assign T97 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign tl_wrap_out = T101 & T98;
  assign T98 = tl_cnt_out == 3'h7;
  assign T144 = reset ? 3'h0 : T99;
  assign T99 = T101 ? T100 : tl_cnt_out;
  assign T100 = tl_cnt_out + 3'h1;
  assign T101 = T103 & is_multibeat;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T102;
  assign T102 = 3'h3 == io_tl_acquire_bits_a_type;
  assign T103 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign io_nasti_w_bits_data = T104;
  assign T104 = io_tl_acquire_bits_data;
  assign io_nasti_w_valid = T105;
  assign T105 = put_valid & aw_ready;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T145 = reset ? 1'h0 : T106;
  assign T106 = T112 ? 1'h0 : T107;
  assign T107 = T108 ? 1'h1 : w_inflight;
  assign T108 = T109 & is_multibeat;
  assign T109 = T111 & T110;
  assign T110 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T111 = w_inflight ^ 1'h1;
  assign T112 = w_inflight & tl_wrap_out;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign io_nasti_aw_bits_user = T113;
  assign T113 = 1'h0;
  assign io_nasti_aw_bits_id = T114;
  assign T114 = T146;
  assign T146 = {1'h0, io_tl_acquire_bits_client_xact_id};
  assign io_nasti_aw_bits_region = T115;
  assign T115 = 4'h0;
  assign io_nasti_aw_bits_qos = T116;
  assign T116 = 4'h0;
  assign io_nasti_aw_bits_prot = T117;
  assign T117 = 3'h0;
  assign io_nasti_aw_bits_cache = T118;
  assign T118 = 4'h0;
  assign io_nasti_aw_bits_lock = T119;
  assign T119 = 1'h0;
  assign io_nasti_aw_bits_burst = T120;
  assign T120 = 2'h1;
  assign io_nasti_aw_bits_size = T121;
  assign T121 = 3'h3;
  assign io_nasti_aw_bits_len = T122;
  assign T122 = T147;
  assign T147 = {5'h0, T123};
  assign T123 = is_multibeat ? 3'h7 : 3'h0;
  assign io_nasti_aw_bits_addr = T124;
  assign T124 = T125;
  assign T125 = {io_tl_acquire_bits_addr_block, T126};
  assign T126 = {io_tl_acquire_bits_addr_beat, T127};
  assign T127 = io_tl_acquire_bits_union[4'hb:4'h9];
  assign io_nasti_aw_valid = T128;
  assign T128 = T130 & T129;
  assign T129 = w_inflight ^ 1'h1;
  assign T130 = put_valid & io_nasti_w_ready;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_acquire_ready = T131;
  assign T131 = has_data ? T133 : T132;
  assign T132 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T133 = aw_ready & io_nasti_w_ready;
  ReorderQueue_1 roq(.clk(clk), .reset(reset),
       .io_enq_ready( roq_io_enq_ready ),
       .io_enq_valid( T37 ),
       .io_enq_bits_data_byteOff( T36 ),
       .io_enq_bits_data_subblock( is_subblock ),
       .io_enq_bits_tag( io_nasti_ar_bits_id ),
       .io_deq_valid( T22 ),
       .io_deq_tag( io_nasti_r_bits_id ),
       .io_deq_data_byteOff( roq_io_deq_data_byteOff ),
       .io_deq_data_subblock( roq_io_deq_data_subblock )
       //.io_deq_matches(  )
  );
  Arbiter_5 gnt_arb(
       .io_in_1_ready( gnt_arb_io_in_1_ready ),
       .io_in_1_valid( io_nasti_b_valid ),
       .io_in_1_bits_addr_beat( T21 ),
       .io_in_1_bits_client_xact_id( T20 ),
       .io_in_1_bits_manager_xact_id( T19 ),
       .io_in_1_bits_is_builtin_type( T18 ),
       .io_in_1_bits_g_type( T17 ),
       .io_in_1_bits_data( T16 ),
       //.io_in_1_bits_client_id(  )
       .io_in_0_ready( gnt_arb_io_in_0_ready ),
       .io_in_0_valid( io_nasti_r_valid ),
       .io_in_0_bits_addr_beat( T8 ),
       .io_in_0_bits_client_xact_id( T7 ),
       .io_in_0_bits_manager_xact_id( T6 ),
       .io_in_0_bits_is_builtin_type( T5 ),
       .io_in_0_bits_g_type( T3 ),
       .io_in_0_bits_data( T0 ),
       //.io_in_0_bits_client_id(  )
       .io_out_ready( io_tl_grant_ready ),
       .io_out_valid( gnt_arb_io_out_valid ),
       .io_out_bits_addr_beat( gnt_arb_io_out_bits_addr_beat ),
       .io_out_bits_client_xact_id( gnt_arb_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( gnt_arb_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( gnt_arb_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( gnt_arb_io_out_bits_g_type ),
       .io_out_bits_data( gnt_arb_io_out_bits_data )
       //.io_out_bits_client_id(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign gnt_arb.io_in_1_bits_client_id = {1{$random}};
    assign gnt_arb.io_in_0_bits_client_id = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else if(T11) begin
      tl_cnt_in <= T10;
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else if(T27) begin
      nasti_cnt_out <= T26;
    end
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else if(T101) begin
      tl_cnt_out <= T100;
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else if(T112) begin
      w_inflight <= 1'h0;
    end else if(T108) begin
      w_inflight <= 1'h1;
    end
  end
endmodule

module ClientTileLinkIOWrapper_1(
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [3:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[3:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[3:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [3:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    //input [25:0] io_out_probe_bits_addr_block
    //input [1:0] io_out_probe_bits_p_type
    input  io_out_release_ready,
    output io_out_release_valid
    //output[1:0] io_out_release_bits_addr_beat
    //output[25:0] io_out_release_bits_addr_block
    //output[3:0] io_out_release_bits_client_xact_id
    //output[2:0] io_out_release_bits_r_type
    //output io_out_release_bits_voluntary
    //output[127:0] io_out_release_bits_data
);



`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_out_release_bits_data = {4{$random}};
//  assign io_out_release_bits_voluntary = {1{$random}};
//  assign io_out_release_bits_r_type = {1{$random}};
//  assign io_out_release_bits_client_xact_id = {1{$random}};
//  assign io_out_release_bits_addr_block = {1{$random}};
//  assign io_out_release_bits_addr_beat = {1{$random}};
// synthesis translate_on
`endif
  assign io_out_release_valid = 1'h0;
  assign io_out_probe_ready = 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_in_grant_bits_data = io_out_grant_bits_data;
  assign io_in_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = io_out_acquire_ready;
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits_data,
    input  io_enq_bits_last,
    input [7:0] io_enq_bits_strb,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits_data,
    output io_deq_bits_last,
    output[7:0] io_deq_bits_strb,
    output io_deq_bits_user,
    output[3:0] io_count
);

  wire[3:0] T0;
  wire[2:0] ptr_diff;
  reg [2:0] R1;
  wire[2:0] T23;
  wire[2:0] T2;
  wire[2:0] T3;
  wire do_deq;
  reg [2:0] R4;
  wire[2:0] T24;
  wire[2:0] T5;
  wire[2:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T25;
  wire T8;
  wire T9;
  wire T10;
  wire[73:0] T11;
  reg [73:0] ram [7:0];
  wire[73:0] T12;
  wire[73:0] T13;
  wire[73:0] T14;
  wire[8:0] T15;
  wire[64:0] T16;
  wire[7:0] T17;
  wire T18;
  wire[63:0] T19;
  wire T20;
  wire empty;
  wire T21;
  wire T22;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T23 = reset ? 3'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 3'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T24 = reset ? 3'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 3'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T25 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T16, T15};
  assign T15 = {io_enq_bits_strb, io_enq_bits_user};
  assign T16 = {io_enq_bits_data, io_enq_bits_last};
  assign io_deq_bits_strb = T17;
  assign T17 = T11[4'h8:1'h1];
  assign io_deq_bits_last = T18;
  assign T18 = T11[4'h9:4'h9];
  assign io_deq_bits_data = T19;
  assign T19 = T11[7'h49:4'ha];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 3'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 3'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_resp,
    input [63:0] io_enq_bits_data,
    input  io_enq_bits_last,
    input [4:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_resp,
    output[63:0] io_deq_bits_data,
    output io_deq_bits_last,
    output[4:0] io_deq_bits_id,
    output io_deq_bits_user,
    output[3:0] io_count
);

  wire[3:0] T0;
  wire[2:0] ptr_diff;
  reg [2:0] R1;
  wire[2:0] T25;
  wire[2:0] T2;
  wire[2:0] T3;
  wire do_deq;
  reg [2:0] R4;
  wire[2:0] T26;
  wire[2:0] T5;
  wire[2:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T27;
  wire T8;
  wire T9;
  wire T10;
  wire[72:0] T11;
  reg [72:0] ram [7:0];
  wire[72:0] T12;
  wire[72:0] T13;
  wire[72:0] T14;
  wire[6:0] T15;
  wire[5:0] T16;
  wire[65:0] T17;
  wire[4:0] T18;
  wire T19;
  wire[63:0] T20;
  wire[1:0] T21;
  wire T22;
  wire empty;
  wire T23;
  wire T24;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T25 = reset ? 3'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 3'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T26 = reset ? 3'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 3'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T27 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T17, T15};
  assign T15 = {io_enq_bits_last, T16};
  assign T16 = {io_enq_bits_id, io_enq_bits_user};
  assign T17 = {io_enq_bits_resp, io_enq_bits_data};
  assign io_deq_bits_id = T18;
  assign T18 = T11[3'h5:1'h1];
  assign io_deq_bits_last = T19;
  assign T19 = T11[3'h6:3'h6];
  assign io_deq_bits_data = T20;
  assign T20 = T11[7'h46:3'h7];
  assign io_deq_bits_resp = T21;
  assign T21 = T11[7'h48:7'h47];
  assign io_deq_valid = T22;
  assign T22 = empty ^ 1'h1;
  assign empty = ptr_match & T23;
  assign T23 = maybe_full ^ 1'h1;
  assign io_enq_ready = T24;
  assign T24 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 3'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 3'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_resp,
    input [4:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_resp,
    output[4:0] io_deq_bits_id,
    output io_deq_bits_user,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire T10;
  wire[7:0] T11;
  reg [7:0] ram [1:0];
  wire[7:0] T12;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[5:0] T15;
  wire[4:0] T16;
  wire[1:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_resp, T15};
  assign T15 = {io_enq_bits_id, io_enq_bits_user};
  assign io_deq_bits_id = T16;
  assign T16 = T11[3'h5:1'h1];
  assign io_deq_bits_resp = T17;
  assign T17 = T11[3'h7:3'h6];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module RTC(input clk, input reset,
    input  io_aw_ready,
    output io_aw_valid,
    output[31:0] io_aw_bits_addr,
    output[7:0] io_aw_bits_len,
    output[2:0] io_aw_bits_size,
    output[1:0] io_aw_bits_burst,
    output io_aw_bits_lock,
    output[3:0] io_aw_bits_cache,
    output[2:0] io_aw_bits_prot,
    output[3:0] io_aw_bits_qos,
    output[3:0] io_aw_bits_region,
    output[4:0] io_aw_bits_id,
    output io_aw_bits_user,
    input  io_w_ready,
    output io_w_valid,
    output[63:0] io_w_bits_data,
    output io_w_bits_last,
    output[7:0] io_w_bits_strb,
    output io_w_bits_user,
    output io_b_ready,
    input  io_b_valid,
    input [1:0] io_b_bits_resp,
    input [4:0] io_b_bits_id,
    input  io_b_bits_user,
    input  io_ar_ready,
    output io_ar_valid,
    //output[31:0] io_ar_bits_addr
    //output[7:0] io_ar_bits_len
    //output[2:0] io_ar_bits_size
    //output[1:0] io_ar_bits_burst
    //output io_ar_bits_lock
    //output[3:0] io_ar_bits_cache
    //output[2:0] io_ar_bits_prot
    //output[3:0] io_ar_bits_qos
    //output[3:0] io_ar_bits_region
    //output[4:0] io_ar_bits_id
    //output io_ar_bits_user
    output io_r_ready,
    input  io_r_valid,
    input [1:0] io_r_bits_resp,
    input [63:0] io_r_bits_data,
    input  io_r_bits_last,
    input [4:0] io_r_bits_id,
    input  io_r_bits_user
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  reg  send_acked_0;
  wire T39;
  wire T3;
  wire T4;
  wire rtc_tick;
  reg [6:0] R5;
  wire[6:0] T40;
  wire[6:0] T6;
  wire[6:0] T7;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire T11;
  wire T41;
  wire T12;
  wire T13;
  wire T14;
  wire[7:0] T15;
  wire T16;
  wire[63:0] T17;
  reg [63:0] rtc;
  wire[63:0] T42;
  wire[63:0] T18;
  wire[63:0] T19;
  reg  sending_data;
  wire T43;
  wire T20;
  wire T21;
  wire[4:0] T22;
  wire[4:0] T44;
  wire coreId;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[2:0] T25;
  wire[3:0] T26;
  wire T27;
  wire[1:0] T28;
  wire[2:0] T29;
  wire[7:0] T30;
  wire[31:0] T31;
  wire[31:0] T45;
  reg [30:0] T32;
  reg  sending_addr;
  wire T46;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    send_acked_0 = {1{$random}};
    R5 = {1{$random}};
    rtc = {2{$random}};
    sending_data = {1{$random}};
    sending_addr = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_ar_bits_user = {1{$random}};
//  assign io_ar_bits_id = {1{$random}};
//  assign io_ar_bits_region = {1{$random}};
//  assign io_ar_bits_qos = {1{$random}};
//  assign io_ar_bits_prot = {1{$random}};
//  assign io_ar_bits_cache = {1{$random}};
//  assign io_ar_bits_lock = {1{$random}};
//  assign io_ar_bits_burst = {1{$random}};
//  assign io_ar_bits_size = {1{$random}};
//  assign io_ar_bits_len = {1{$random}};
//  assign io_ar_bits_addr = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T13 | send_acked_0;
  assign T39 = reset ? 1'h1 : T3;
  assign T3 = T8 ? 1'h1 : T4;
  assign T4 = rtc_tick ? 1'h0 : send_acked_0;
  assign rtc_tick = R5 == 7'h63;
  assign T40 = reset ? 7'h0 : T6;
  assign T6 = rtc_tick ? 7'h0 : T7;
  assign T7 = R5 + 7'h1;
  assign T8 = T12 & T9;
  assign T9 = T10[1'h0:1'h0];
  assign T10 = 1'h1 << T11;
  assign T11 = T41;
  assign T41 = io_b_bits_id[1'h0:1'h0];
  assign T12 = io_b_ready & io_b_valid;
  assign T13 = rtc_tick ^ 1'h1;
  assign io_r_ready = 1'h0;
  assign io_ar_valid = 1'h0;
  assign io_b_ready = 1'h1;
  assign io_w_bits_user = T14;
  assign T14 = 1'h0;
  assign io_w_bits_strb = T15;
  assign T15 = 8'hff;
  assign io_w_bits_last = T16;
  assign T16 = 1'h1;
  assign io_w_bits_data = T17;
  assign T17 = rtc;
  assign T42 = reset ? 64'h0 : T18;
  assign T18 = rtc_tick ? T19 : rtc;
  assign T19 = rtc + 64'h1;
  assign io_w_valid = sending_data;
  assign T43 = reset ? 1'h0 : T20;
  assign T20 = rtc_tick ? 1'h1 : sending_data;
  assign io_aw_bits_user = T21;
  assign T21 = 1'h0;
  assign io_aw_bits_id = T22;
  assign T22 = T44;
  assign T44 = {4'h0, coreId};
  assign coreId = 1'h0;
  assign io_aw_bits_region = T23;
  assign T23 = 4'h0;
  assign io_aw_bits_qos = T24;
  assign T24 = 4'h0;
  assign io_aw_bits_prot = T25;
  assign T25 = 3'h0;
  assign io_aw_bits_cache = T26;
  assign T26 = 4'h0;
  assign io_aw_bits_lock = T27;
  assign T27 = 1'h0;
  assign io_aw_bits_burst = T28;
  assign T28 = 2'h1;
  assign io_aw_bits_size = T29;
  assign T29 = 3'h3;
  assign io_aw_bits_len = T30;
  assign T30 = 8'h0;
  assign io_aw_bits_addr = T31;
  assign T31 = T45;
  assign T45 = {1'h0, T32};
  always @(*) case (coreId)
    0: T32 = 31'h40003808;
    default: begin
      T32 = 31'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T32 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign io_aw_valid = sending_addr;
  assign T46 = reset ? 1'h0 : T34;
  assign T34 = T38 ? 1'h0 : T35;
  assign T35 = T37 ? 1'h0 : T36;
  assign T36 = rtc_tick ? 1'h1 : sending_addr;
  assign T37 = io_aw_ready & io_aw_valid;
  assign T38 = io_w_ready & io_w_valid;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Not all clocks were updated for rtc tick");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      send_acked_0 <= 1'h1;
    end else if(T8) begin
      send_acked_0 <= 1'h1;
    end else if(rtc_tick) begin
      send_acked_0 <= 1'h0;
    end
    if(reset) begin
      R5 <= 7'h0;
    end else if(rtc_tick) begin
      R5 <= 7'h0;
    end else begin
      R5 <= T7;
    end
    if(reset) begin
      rtc <= 64'h0;
    end else if(rtc_tick) begin
      rtc <= T19;
    end
    if(reset) begin
      sending_data <= 1'h0;
    end else if(rtc_tick) begin
      sending_data <= 1'h1;
    end
    if(reset) begin
      sending_addr <= 1'h0;
    end else if(T38) begin
      sending_addr <= 1'h0;
    end else if(T37) begin
      sending_addr <= 1'h0;
    end else if(rtc_tick) begin
      sending_addr <= 1'h1;
    end
  end
endmodule

module SMIIONastiReadIOConverter_0(input clk, input reset,
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [4:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[4:0] io_r_bits_id,
    output io_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[11:0] io_smi_req_bits_addr,
    //output[63:0] io_smi_req_bits_data
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire T0;
  reg [1:0] state;
  wire[1:0] T60;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  reg  nWords;
  wire T61;
  wire[7:0] T7;
  wire[7:0] T62;
  wire T8;
  wire T9;
  wire T10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg  recvInd;
  wire T63;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire T21;
  reg [11:0] addr;
  wire[11:0] T22;
  wire[11:0] T23;
  wire[11:0] T24;
  wire[11:0] T25;
  wire T26;
  wire T27;
  wire T28;
  reg  sendDone;
  wire T64;
  wire T29;
  wire T30;
  wire T31;
  reg  sendInd;
  wire T65;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[4:0] T37;
  reg [4:0] id;
  wire[4:0] T38;
  wire T39;
  wire T40;
  reg [7:0] nBeats;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[63:0] T44;
  wire[63:0] T45;
  reg [63:0] buffer_0;
  wire[63:0] T66;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[5:0] T49;
  reg [2:0] byteOff;
  wire[2:0] T50;
  wire[2:0] T51;
  wire[2:0] T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    nWords = {1{$random}};
    recvInd = {1{$random}};
    addr = {1{$random}};
    sendDone = {1{$random}};
    sendInd = {1{$random}};
    id = {1{$random}};
    nBeats = {1{$random}};
    buffer_0 = {2{$random}};
    byteOff = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_smi_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
  assign io_smi_resp_ready = T0;
  assign T0 = state == 2'h1;
  assign T60 = reset ? 2'h0 : T1;
  assign T1 = T21 ? T20 : T2;
  assign T2 = T5 ? 2'h2 : T3;
  assign T3 = T4 ? 2'h1 : state;
  assign T4 = io_ar_ready & io_ar_valid;
  assign T5 = T19 & T6;
  assign T6 = recvInd == nWords;
  assign T61 = T7[1'h0:1'h0];
  assign T7 = T14 ? T11 : T62;
  assign T62 = {7'h0, T8};
  assign T8 = T9 ? 1'h0 : nWords;
  assign T9 = T4 & T10;
  assign T10 = io_ar_bits_size < 3'h3;
  assign T11 = T12 - 8'h1;
  assign T12 = 1'h1 << T13;
  assign T13 = io_ar_bits_size - 3'h3;
  assign T14 = T4 & T15;
  assign T15 = T10 ^ 1'h1;
  assign T63 = reset ? 1'h0 : T16;
  assign T16 = T21 ? 1'h0 : T17;
  assign T17 = T19 ? T18 : recvInd;
  assign T18 = recvInd + 1'h1;
  assign T19 = io_smi_resp_ready & io_smi_resp_valid;
  assign T20 = io_r_bits_last ? 2'h0 : 2'h1;
  assign T21 = io_r_ready & io_r_valid;
  assign io_smi_req_bits_addr = addr;
  assign T22 = T26 ? T25 : T23;
  assign T23 = T4 ? T24 : addr;
  assign T24 = io_ar_bits_addr[4'he:2'h3];
  assign T25 = addr + 12'h1;
  assign T26 = io_smi_req_ready & io_smi_req_valid;
  assign io_smi_req_bits_rw = 1'h0;
  assign io_smi_req_valid = T27;
  assign T27 = T35 & T28;
  assign T28 = sendDone ^ 1'h1;
  assign T64 = reset ? 1'h0 : T29;
  assign T29 = T21 ? 1'h0 : T30;
  assign T30 = T26 ? T31 : sendDone;
  assign T31 = sendInd == nWords;
  assign T65 = reset ? 1'h0 : T32;
  assign T32 = T21 ? 1'h0 : T33;
  assign T33 = T26 ? T34 : sendInd;
  assign T34 = sendInd + 1'h1;
  assign T35 = state == 2'h1;
  assign io_r_bits_user = T36;
  assign T36 = 1'h0;
  assign io_r_bits_id = T37;
  assign T37 = id;
  assign T38 = T4 ? io_ar_bits_id : id;
  assign io_r_bits_last = T39;
  assign T39 = T40;
  assign T40 = nBeats == 8'h0;
  assign T41 = T21 ? T43 : T42;
  assign T42 = T4 ? io_ar_bits_len : nBeats;
  assign T43 = nBeats - 8'h1;
  assign io_r_bits_data = T44;
  assign T44 = T45;
  assign T45 = buffer_0;
  assign T66 = reset ? 64'h0 : T46;
  assign T46 = T21 ? 64'h0 : T47;
  assign T47 = T53 ? T48 : buffer_0;
  assign T48 = io_smi_resp_bits >> T49;
  assign T49 = {byteOff, 3'h0};
  assign T50 = T14 ? 3'h0 : T51;
  assign T51 = T9 ? T52 : byteOff;
  assign T52 = io_ar_bits_addr[2'h2:1'h0];
  assign T53 = T19 & T54;
  assign T54 = T55[1'h0:1'h0];
  assign T55 = 1'h1 << T56;
  assign T56 = recvInd;
  assign io_r_bits_resp = T57;
  assign T57 = 2'h0;
  assign io_r_valid = T58;
  assign T58 = state == 2'h2;
  assign io_ar_ready = T59;
  assign T59 = state == 2'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T21) begin
      state <= T20;
    end else if(T5) begin
      state <= 2'h2;
    end else if(T4) begin
      state <= 2'h1;
    end
    nWords <= T61;
    if(reset) begin
      recvInd <= 1'h0;
    end else if(T21) begin
      recvInd <= 1'h0;
    end else if(T19) begin
      recvInd <= T18;
    end
    if(T26) begin
      addr <= T25;
    end else if(T4) begin
      addr <= T24;
    end
    if(reset) begin
      sendDone <= 1'h0;
    end else if(T21) begin
      sendDone <= 1'h0;
    end else if(T26) begin
      sendDone <= T31;
    end
    if(reset) begin
      sendInd <= 1'h0;
    end else if(T21) begin
      sendInd <= 1'h0;
    end else if(T26) begin
      sendInd <= T34;
    end
    if(T4) begin
      id <= io_ar_bits_id;
    end
    if(T21) begin
      nBeats <= T43;
    end else if(T4) begin
      nBeats <= io_ar_bits_len;
    end
    if(reset) begin
      buffer_0 <= 64'h0;
    end else if(T21) begin
      buffer_0 <= 64'h0;
    end else if(T53) begin
      buffer_0 <= T48;
    end
    if(T14) begin
      byteOff <= 3'h0;
    end else if(T9) begin
      byteOff <= T52;
    end
  end
endmodule

module SMIIONastiWriteIOConverter_0(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [4:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    output[1:0] io_b_bits_resp,
    output[4:0] io_b_bits_id,
    output io_b_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[11:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  reg [2:0] state;
  wire[2:0] T52;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire[2:0] T13;
  reg  last;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  strb;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[255:0] T22;
  wire[255:0] T53;
  wire[255:0] T23;
  wire[255:0] T24;
  wire[7:0] T25;
  reg [2:0] size;
  wire[2:0] T26;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg [63:0] data;
  wire[63:0] T36;
  wire[63:0] T37;
  reg [11:0] addr;
  wire[11:0] T39;
  wire[11:0] T40;
  wire[11:0] T41;
  wire[11:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[4:0] T46;
  reg [4:0] id;
  wire[4:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire T51;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    last = {1{$random}};
    strb = {1{$random}};
    size = {1{$random}};
    data = {2{$random}};
    addr = {1{$random}};
    id = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T4 | T3;
  assign T3 = 3'h3 <= io_aw_bits_size;
  assign T4 = io_aw_valid ^ 1'h1;
  assign io_smi_resp_ready = T5;
  assign T5 = state == 3'h3;
  assign T52 = reset ? 3'h0 : T6;
  assign T6 = T35 ? 3'h0 : T7;
  assign T7 = T34 ? 3'h4 : T8;
  assign T8 = T16 ? T13 : T9;
  assign T9 = T12 ? 3'h2 : T10;
  assign T10 = T11 ? 3'h1 : state;
  assign T11 = io_aw_ready & io_aw_valid;
  assign T12 = io_w_ready & io_w_valid;
  assign T13 = last ? 3'h3 : 3'h1;
  assign T14 = T12 ? io_w_bits_last : T15;
  assign T15 = T11 ? 1'h0 : last;
  assign T16 = T33 & T17;
  assign T17 = strb == 1'h0;
  assign T18 = T28 ? 1'h0 : T19;
  assign T19 = T12 ? T20 : strb;
  assign T20 = T21;
  assign T21 = T22[1'h0:1'h0];
  assign T22 = T23 & T53;
  assign T53 = {248'h0, io_w_bits_strb};
  assign T23 = T24 - 256'h1;
  assign T24 = 1'h1 << T25;
  assign T25 = 1'h1 << size;
  assign T26 = T11 ? io_aw_bits_size : size;
  assign T28 = T33 & T29;
  assign T29 = T32 & T30;
  assign T30 = io_smi_req_ready | T31;
  assign T31 = strb ^ 1'h1;
  assign T32 = T17 ^ 1'h1;
  assign T33 = state == 3'h2;
  assign T34 = io_smi_resp_ready & io_smi_resp_valid;
  assign T35 = io_b_ready & io_b_valid;
  assign io_smi_req_bits_data = data;
  assign T36 = T28 ? 64'h0 : T37;
  assign T37 = T12 ? io_w_bits_data : data;
  assign io_smi_req_bits_addr = addr;
  assign T39 = T28 ? T42 : T40;
  assign T40 = T11 ? T41 : addr;
  assign T41 = io_aw_bits_addr[4'he:2'h3];
  assign T42 = addr + 12'h1;
  assign io_smi_req_bits_rw = 1'h1;
  assign io_smi_req_valid = T43;
  assign T43 = T44 & strb;
  assign T44 = state == 3'h2;
  assign io_b_bits_user = T45;
  assign T45 = 1'h0;
  assign io_b_bits_id = T46;
  assign T46 = id;
  assign T47 = T11 ? io_aw_bits_id : id;
  assign io_b_bits_resp = T48;
  assign T48 = 2'h0;
  assign io_b_valid = T49;
  assign T49 = state == 3'h4;
  assign io_w_ready = T50;
  assign T50 = state == 3'h1;
  assign io_aw_ready = T51;
  assign T51 = state == 3'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Nasti size must be >= SMI size");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h4;
    end else if(T16) begin
      state <= T13;
    end else if(T12) begin
      state <= 3'h2;
    end else if(T11) begin
      state <= 3'h1;
    end
    if(T12) begin
      last <= io_w_bits_last;
    end else if(T11) begin
      last <= 1'h0;
    end
    if(T28) begin
      strb <= 1'h0;
    end else if(T12) begin
      strb <= T20;
    end
    if(T11) begin
      size <= io_aw_bits_size;
    end
    if(T28) begin
      data <= 64'h0;
    end else if(T12) begin
      data <= io_w_bits_data;
    end
    if(T28) begin
      addr <= T42;
    end else if(T11) begin
      addr <= T41;
    end
    if(T11) begin
      id <= io_aw_bits_id;
    end
  end
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_rw,
    input [11:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_rw,
    input [11:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_rw,
    output[11:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T27;
  wire T3;
  wire T4;
  wire[63:0] T5;
  wire T6;
  wire[11:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T27 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_data = T5;
  assign T5 = T6 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T6 = chosen;
  assign io_out_bits_addr = T7;
  assign T7 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_rw = T8;
  assign T8 = T6 ? io_in_1_bits_rw : io_in_0_bits_rw;
  assign io_out_valid = T9;
  assign T9 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = T18 | T12;
  assign T12 = T13 ^ 1'h1;
  assign T13 = T16 | T14;
  assign T14 = io_in_1_valid & T15;
  assign T15 = last_grant < 1'h1;
  assign T16 = io_in_0_valid & T17;
  assign T17 = last_grant < 1'h0;
  assign T18 = last_grant < 1'h0;
  assign io_in_1_ready = T19;
  assign T19 = T20 & io_out_ready;
  assign T20 = T24 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = T23 | io_in_0_valid;
  assign T23 = T16 | T14;
  assign T24 = T26 & T25;
  assign T25 = last_grant < 1'h1;
  assign T26 = T16 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module SMIArbiter_0(input clk, input reset,
    output io_in_1_req_ready,
    input  io_in_1_req_valid,
    input  io_in_1_req_bits_rw,
    input [11:0] io_in_1_req_bits_addr,
    input [63:0] io_in_1_req_bits_data,
    input  io_in_1_resp_ready,
    output io_in_1_resp_valid,
    output[63:0] io_in_1_resp_bits,
    output io_in_0_req_ready,
    input  io_in_0_req_valid,
    input  io_in_0_req_bits_rw,
    input [11:0] io_in_0_req_bits_addr,
    input [63:0] io_in_0_req_bits_data,
    input  io_in_0_resp_ready,
    output io_in_0_resp_valid,
    output[63:0] io_in_0_resp_bits,
    input  io_out_req_ready,
    output io_out_req_valid,
    output io_out_req_bits_rw,
    output[11:0] io_out_req_bits_addr,
    output[63:0] io_out_req_bits_data,
    output io_out_resp_ready,
    input  io_out_resp_valid,
    input [63:0] io_out_resp_bits
);

  wire T0;
  wire T1;
  reg  wait_resp;
  wire T15;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  choice;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire req_arb_io_in_1_ready;
  wire req_arb_io_in_0_ready;
  wire req_arb_io_out_valid;
  wire req_arb_io_out_bits_rw;
  wire[11:0] req_arb_io_out_bits_addr;
  wire[63:0] req_arb_io_out_bits_data;
  wire req_arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wait_resp = {1{$random}};
    choice = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_out_req_ready & T1;
  assign T1 = wait_resp ^ 1'h1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = T5 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : wait_resp;
  assign T4 = io_out_req_ready & io_out_req_valid;
  assign T5 = io_out_resp_ready & io_out_resp_valid;
  assign io_out_resp_ready = T6;
  assign T6 = T7 ? io_in_1_resp_ready : io_in_0_resp_ready;
  assign T7 = choice;
  assign T8 = T4 ? req_arb_io_chosen : choice;
  assign io_out_req_bits_data = req_arb_io_out_bits_data;
  assign io_out_req_bits_addr = req_arb_io_out_bits_addr;
  assign io_out_req_bits_rw = req_arb_io_out_bits_rw;
  assign io_out_req_valid = T9;
  assign T9 = req_arb_io_out_valid & T10;
  assign T10 = wait_resp ^ 1'h1;
  assign io_in_0_resp_bits = io_out_resp_bits;
  assign io_in_0_resp_valid = T11;
  assign T11 = io_out_resp_valid & T12;
  assign T12 = choice == 1'h0;
  assign io_in_0_req_ready = req_arb_io_in_0_ready;
  assign io_in_1_resp_bits = io_out_resp_bits;
  assign io_in_1_resp_valid = T13;
  assign T13 = io_out_resp_valid & T14;
  assign T14 = choice == 1'h1;
  assign io_in_1_req_ready = req_arb_io_in_1_ready;
  RRArbiter_0 req_arb(.clk(clk), .reset(reset),
       .io_in_1_ready( req_arb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_req_valid ),
       .io_in_1_bits_rw( io_in_1_req_bits_rw ),
       .io_in_1_bits_addr( io_in_1_req_bits_addr ),
       .io_in_1_bits_data( io_in_1_req_bits_data ),
       .io_in_0_ready( req_arb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_req_valid ),
       .io_in_0_bits_rw( io_in_0_req_bits_rw ),
       .io_in_0_bits_addr( io_in_0_req_bits_addr ),
       .io_in_0_bits_data( io_in_0_req_bits_data ),
       .io_out_ready( T0 ),
       .io_out_valid( req_arb_io_out_valid ),
       .io_out_bits_rw( req_arb_io_out_bits_rw ),
       .io_out_bits_addr( req_arb_io_out_bits_addr ),
       .io_out_bits_data( req_arb_io_out_bits_data ),
       .io_chosen( req_arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      wait_resp <= 1'h0;
    end else if(T5) begin
      wait_resp <= 1'h0;
    end else if(T4) begin
      wait_resp <= 1'h1;
    end
    if(T4) begin
      choice <= req_arb_io_chosen;
    end
  end
endmodule

module SMIIONastiIOConverter_0(input clk, input reset,
    output io_nasti_aw_ready,
    input  io_nasti_aw_valid,
    input [31:0] io_nasti_aw_bits_addr,
    input [7:0] io_nasti_aw_bits_len,
    input [2:0] io_nasti_aw_bits_size,
    input [1:0] io_nasti_aw_bits_burst,
    input  io_nasti_aw_bits_lock,
    input [3:0] io_nasti_aw_bits_cache,
    input [2:0] io_nasti_aw_bits_prot,
    input [3:0] io_nasti_aw_bits_qos,
    input [3:0] io_nasti_aw_bits_region,
    input [4:0] io_nasti_aw_bits_id,
    input  io_nasti_aw_bits_user,
    output io_nasti_w_ready,
    input  io_nasti_w_valid,
    input [63:0] io_nasti_w_bits_data,
    input  io_nasti_w_bits_last,
    input [7:0] io_nasti_w_bits_strb,
    input  io_nasti_w_bits_user,
    input  io_nasti_b_ready,
    output io_nasti_b_valid,
    output[1:0] io_nasti_b_bits_resp,
    output[4:0] io_nasti_b_bits_id,
    output io_nasti_b_bits_user,
    output io_nasti_ar_ready,
    input  io_nasti_ar_valid,
    input [31:0] io_nasti_ar_bits_addr,
    input [7:0] io_nasti_ar_bits_len,
    input [2:0] io_nasti_ar_bits_size,
    input [1:0] io_nasti_ar_bits_burst,
    input  io_nasti_ar_bits_lock,
    input [3:0] io_nasti_ar_bits_cache,
    input [2:0] io_nasti_ar_bits_prot,
    input [3:0] io_nasti_ar_bits_qos,
    input [3:0] io_nasti_ar_bits_region,
    input [4:0] io_nasti_ar_bits_id,
    input  io_nasti_ar_bits_user,
    input  io_nasti_r_ready,
    output io_nasti_r_valid,
    output[1:0] io_nasti_r_bits_resp,
    output[63:0] io_nasti_r_bits_data,
    output io_nasti_r_bits_last,
    output[4:0] io_nasti_r_bits_id,
    output io_nasti_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[11:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire reader_io_ar_ready;
  wire reader_io_r_valid;
  wire[1:0] reader_io_r_bits_resp;
  wire[63:0] reader_io_r_bits_data;
  wire reader_io_r_bits_last;
  wire[4:0] reader_io_r_bits_id;
  wire reader_io_r_bits_user;
  wire reader_io_smi_req_valid;
  wire reader_io_smi_req_bits_rw;
  wire[11:0] reader_io_smi_req_bits_addr;
  wire reader_io_smi_resp_ready;
  wire writer_io_aw_ready;
  wire writer_io_w_ready;
  wire writer_io_b_valid;
  wire[1:0] writer_io_b_bits_resp;
  wire[4:0] writer_io_b_bits_id;
  wire writer_io_b_bits_user;
  wire writer_io_smi_req_valid;
  wire writer_io_smi_req_bits_rw;
  wire[11:0] writer_io_smi_req_bits_addr;
  wire[63:0] writer_io_smi_req_bits_data;
  wire writer_io_smi_resp_ready;
  wire arb_io_in_1_req_ready;
  wire arb_io_in_1_resp_valid;
  wire[63:0] arb_io_in_1_resp_bits;
  wire arb_io_in_0_req_ready;
  wire arb_io_in_0_resp_valid;
  wire[63:0] arb_io_in_0_resp_bits;
  wire arb_io_out_req_valid;
  wire arb_io_out_req_bits_rw;
  wire[11:0] arb_io_out_req_bits_addr;
  wire[63:0] arb_io_out_req_bits_data;
  wire arb_io_out_resp_ready;


  assign io_smi_resp_ready = arb_io_out_resp_ready;
  assign io_smi_req_bits_data = arb_io_out_req_bits_data;
  assign io_smi_req_bits_addr = arb_io_out_req_bits_addr;
  assign io_smi_req_bits_rw = arb_io_out_req_bits_rw;
  assign io_smi_req_valid = arb_io_out_req_valid;
  assign io_nasti_r_bits_user = reader_io_r_bits_user;
  assign io_nasti_r_bits_id = reader_io_r_bits_id;
  assign io_nasti_r_bits_last = reader_io_r_bits_last;
  assign io_nasti_r_bits_data = reader_io_r_bits_data;
  assign io_nasti_r_bits_resp = reader_io_r_bits_resp;
  assign io_nasti_r_valid = reader_io_r_valid;
  assign io_nasti_ar_ready = reader_io_ar_ready;
  assign io_nasti_b_bits_user = writer_io_b_bits_user;
  assign io_nasti_b_bits_id = writer_io_b_bits_id;
  assign io_nasti_b_bits_resp = writer_io_b_bits_resp;
  assign io_nasti_b_valid = writer_io_b_valid;
  assign io_nasti_w_ready = writer_io_w_ready;
  assign io_nasti_aw_ready = writer_io_aw_ready;
  SMIIONastiReadIOConverter_0 reader(.clk(clk), .reset(reset),
       .io_ar_ready( reader_io_ar_ready ),
       .io_ar_valid( io_nasti_ar_valid ),
       .io_ar_bits_addr( io_nasti_ar_bits_addr ),
       .io_ar_bits_len( io_nasti_ar_bits_len ),
       .io_ar_bits_size( io_nasti_ar_bits_size ),
       .io_ar_bits_burst( io_nasti_ar_bits_burst ),
       .io_ar_bits_lock( io_nasti_ar_bits_lock ),
       .io_ar_bits_cache( io_nasti_ar_bits_cache ),
       .io_ar_bits_prot( io_nasti_ar_bits_prot ),
       .io_ar_bits_qos( io_nasti_ar_bits_qos ),
       .io_ar_bits_region( io_nasti_ar_bits_region ),
       .io_ar_bits_id( io_nasti_ar_bits_id ),
       .io_ar_bits_user( io_nasti_ar_bits_user ),
       .io_r_ready( io_nasti_r_ready ),
       .io_r_valid( reader_io_r_valid ),
       .io_r_bits_resp( reader_io_r_bits_resp ),
       .io_r_bits_data( reader_io_r_bits_data ),
       .io_r_bits_last( reader_io_r_bits_last ),
       .io_r_bits_id( reader_io_r_bits_id ),
       .io_r_bits_user( reader_io_r_bits_user ),
       .io_smi_req_ready( arb_io_in_0_req_ready ),
       .io_smi_req_valid( reader_io_smi_req_valid ),
       .io_smi_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_smi_req_bits_data(  )
       .io_smi_resp_ready( reader_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_0_resp_valid ),
       .io_smi_resp_bits( arb_io_in_0_resp_bits )
  );
  SMIIONastiWriteIOConverter_0 writer(.clk(clk), .reset(reset),
       .io_aw_ready( writer_io_aw_ready ),
       .io_aw_valid( io_nasti_aw_valid ),
       .io_aw_bits_addr( io_nasti_aw_bits_addr ),
       .io_aw_bits_len( io_nasti_aw_bits_len ),
       .io_aw_bits_size( io_nasti_aw_bits_size ),
       .io_aw_bits_burst( io_nasti_aw_bits_burst ),
       .io_aw_bits_lock( io_nasti_aw_bits_lock ),
       .io_aw_bits_cache( io_nasti_aw_bits_cache ),
       .io_aw_bits_prot( io_nasti_aw_bits_prot ),
       .io_aw_bits_qos( io_nasti_aw_bits_qos ),
       .io_aw_bits_region( io_nasti_aw_bits_region ),
       .io_aw_bits_id( io_nasti_aw_bits_id ),
       .io_aw_bits_user( io_nasti_aw_bits_user ),
       .io_w_ready( writer_io_w_ready ),
       .io_w_valid( io_nasti_w_valid ),
       .io_w_bits_data( io_nasti_w_bits_data ),
       .io_w_bits_last( io_nasti_w_bits_last ),
       .io_w_bits_strb( io_nasti_w_bits_strb ),
       .io_w_bits_user( io_nasti_w_bits_user ),
       .io_b_ready( io_nasti_b_ready ),
       .io_b_valid( writer_io_b_valid ),
       .io_b_bits_resp( writer_io_b_bits_resp ),
       .io_b_bits_id( writer_io_b_bits_id ),
       .io_b_bits_user( writer_io_b_bits_user ),
       .io_smi_req_ready( arb_io_in_1_req_ready ),
       .io_smi_req_valid( writer_io_smi_req_valid ),
       .io_smi_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( writer_io_smi_req_bits_data ),
       .io_smi_resp_ready( writer_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_1_resp_valid ),
       .io_smi_resp_bits( arb_io_in_1_resp_bits )
  );
  SMIArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_1_req_ready( arb_io_in_1_req_ready ),
       .io_in_1_req_valid( writer_io_smi_req_valid ),
       .io_in_1_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_in_1_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_in_1_req_bits_data( writer_io_smi_req_bits_data ),
       .io_in_1_resp_ready( writer_io_smi_resp_ready ),
       .io_in_1_resp_valid( arb_io_in_1_resp_valid ),
       .io_in_1_resp_bits( arb_io_in_1_resp_bits ),
       .io_in_0_req_ready( arb_io_in_0_req_ready ),
       .io_in_0_req_valid( reader_io_smi_req_valid ),
       .io_in_0_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_in_0_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_in_0_req_bits_data(  )
       .io_in_0_resp_ready( reader_io_smi_resp_ready ),
       .io_in_0_resp_valid( arb_io_in_0_resp_valid ),
       .io_in_0_resp_bits( arb_io_in_0_resp_bits ),
       .io_out_req_ready( io_smi_req_ready ),
       .io_out_req_valid( arb_io_out_req_valid ),
       .io_out_req_bits_rw( arb_io_out_req_bits_rw ),
       .io_out_req_bits_addr( arb_io_out_req_bits_addr ),
       .io_out_req_bits_data( arb_io_out_req_bits_data ),
       .io_out_resp_ready( arb_io_out_resp_ready ),
       .io_out_resp_valid( io_smi_resp_valid ),
       .io_out_resp_bits( io_smi_resp_bits )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign arb.io_in_0_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
endmodule

module SMIIONastiReadIOConverter_1(input clk, input reset,
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [4:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[4:0] io_r_bits_id,
    output io_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[5:0] io_smi_req_bits_addr,
    //output[63:0] io_smi_req_bits_data
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire T0;
  reg [1:0] state;
  wire[1:0] T60;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  reg  nWords;
  wire T61;
  wire[7:0] T7;
  wire[7:0] T62;
  wire T8;
  wire T9;
  wire T10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg  recvInd;
  wire T63;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire T21;
  reg [5:0] addr;
  wire[5:0] T22;
  wire[5:0] T23;
  wire[5:0] T24;
  wire[5:0] T25;
  wire T26;
  wire T27;
  wire T28;
  reg  sendDone;
  wire T64;
  wire T29;
  wire T30;
  wire T31;
  reg  sendInd;
  wire T65;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[4:0] T37;
  reg [4:0] id;
  wire[4:0] T38;
  wire T39;
  wire T40;
  reg [7:0] nBeats;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[63:0] T44;
  wire[63:0] T45;
  reg [63:0] buffer_0;
  wire[63:0] T66;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[5:0] T49;
  reg [2:0] byteOff;
  wire[2:0] T50;
  wire[2:0] T51;
  wire[2:0] T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    nWords = {1{$random}};
    recvInd = {1{$random}};
    addr = {1{$random}};
    sendDone = {1{$random}};
    sendInd = {1{$random}};
    id = {1{$random}};
    nBeats = {1{$random}};
    buffer_0 = {2{$random}};
    byteOff = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_smi_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
  assign io_smi_resp_ready = T0;
  assign T0 = state == 2'h1;
  assign T60 = reset ? 2'h0 : T1;
  assign T1 = T21 ? T20 : T2;
  assign T2 = T5 ? 2'h2 : T3;
  assign T3 = T4 ? 2'h1 : state;
  assign T4 = io_ar_ready & io_ar_valid;
  assign T5 = T19 & T6;
  assign T6 = recvInd == nWords;
  assign T61 = T7[1'h0:1'h0];
  assign T7 = T14 ? T11 : T62;
  assign T62 = {7'h0, T8};
  assign T8 = T9 ? 1'h0 : nWords;
  assign T9 = T4 & T10;
  assign T10 = io_ar_bits_size < 3'h3;
  assign T11 = T12 - 8'h1;
  assign T12 = 1'h1 << T13;
  assign T13 = io_ar_bits_size - 3'h3;
  assign T14 = T4 & T15;
  assign T15 = T10 ^ 1'h1;
  assign T63 = reset ? 1'h0 : T16;
  assign T16 = T21 ? 1'h0 : T17;
  assign T17 = T19 ? T18 : recvInd;
  assign T18 = recvInd + 1'h1;
  assign T19 = io_smi_resp_ready & io_smi_resp_valid;
  assign T20 = io_r_bits_last ? 2'h0 : 2'h1;
  assign T21 = io_r_ready & io_r_valid;
  assign io_smi_req_bits_addr = addr;
  assign T22 = T26 ? T25 : T23;
  assign T23 = T4 ? T24 : addr;
  assign T24 = io_ar_bits_addr[4'h8:2'h3];
  assign T25 = addr + 6'h1;
  assign T26 = io_smi_req_ready & io_smi_req_valid;
  assign io_smi_req_bits_rw = 1'h0;
  assign io_smi_req_valid = T27;
  assign T27 = T35 & T28;
  assign T28 = sendDone ^ 1'h1;
  assign T64 = reset ? 1'h0 : T29;
  assign T29 = T21 ? 1'h0 : T30;
  assign T30 = T26 ? T31 : sendDone;
  assign T31 = sendInd == nWords;
  assign T65 = reset ? 1'h0 : T32;
  assign T32 = T21 ? 1'h0 : T33;
  assign T33 = T26 ? T34 : sendInd;
  assign T34 = sendInd + 1'h1;
  assign T35 = state == 2'h1;
  assign io_r_bits_user = T36;
  assign T36 = 1'h0;
  assign io_r_bits_id = T37;
  assign T37 = id;
  assign T38 = T4 ? io_ar_bits_id : id;
  assign io_r_bits_last = T39;
  assign T39 = T40;
  assign T40 = nBeats == 8'h0;
  assign T41 = T21 ? T43 : T42;
  assign T42 = T4 ? io_ar_bits_len : nBeats;
  assign T43 = nBeats - 8'h1;
  assign io_r_bits_data = T44;
  assign T44 = T45;
  assign T45 = buffer_0;
  assign T66 = reset ? 64'h0 : T46;
  assign T46 = T21 ? 64'h0 : T47;
  assign T47 = T53 ? T48 : buffer_0;
  assign T48 = io_smi_resp_bits >> T49;
  assign T49 = {byteOff, 3'h0};
  assign T50 = T14 ? 3'h0 : T51;
  assign T51 = T9 ? T52 : byteOff;
  assign T52 = io_ar_bits_addr[2'h2:1'h0];
  assign T53 = T19 & T54;
  assign T54 = T55[1'h0:1'h0];
  assign T55 = 1'h1 << T56;
  assign T56 = recvInd;
  assign io_r_bits_resp = T57;
  assign T57 = 2'h0;
  assign io_r_valid = T58;
  assign T58 = state == 2'h2;
  assign io_ar_ready = T59;
  assign T59 = state == 2'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T21) begin
      state <= T20;
    end else if(T5) begin
      state <= 2'h2;
    end else if(T4) begin
      state <= 2'h1;
    end
    nWords <= T61;
    if(reset) begin
      recvInd <= 1'h0;
    end else if(T21) begin
      recvInd <= 1'h0;
    end else if(T19) begin
      recvInd <= T18;
    end
    if(T26) begin
      addr <= T25;
    end else if(T4) begin
      addr <= T24;
    end
    if(reset) begin
      sendDone <= 1'h0;
    end else if(T21) begin
      sendDone <= 1'h0;
    end else if(T26) begin
      sendDone <= T31;
    end
    if(reset) begin
      sendInd <= 1'h0;
    end else if(T21) begin
      sendInd <= 1'h0;
    end else if(T26) begin
      sendInd <= T34;
    end
    if(T4) begin
      id <= io_ar_bits_id;
    end
    if(T21) begin
      nBeats <= T43;
    end else if(T4) begin
      nBeats <= io_ar_bits_len;
    end
    if(reset) begin
      buffer_0 <= 64'h0;
    end else if(T21) begin
      buffer_0 <= 64'h0;
    end else if(T53) begin
      buffer_0 <= T48;
    end
    if(T14) begin
      byteOff <= 3'h0;
    end else if(T9) begin
      byteOff <= T52;
    end
  end
endmodule

module SMIIONastiWriteIOConverter_1(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [4:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    output[1:0] io_b_bits_resp,
    output[4:0] io_b_bits_id,
    output io_b_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[5:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  reg [2:0] state;
  wire[2:0] T52;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire[2:0] T13;
  reg  last;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  strb;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[255:0] T22;
  wire[255:0] T53;
  wire[255:0] T23;
  wire[255:0] T24;
  wire[7:0] T25;
  reg [2:0] size;
  wire[2:0] T26;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg [63:0] data;
  wire[63:0] T36;
  wire[63:0] T37;
  reg [5:0] addr;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[4:0] T46;
  reg [4:0] id;
  wire[4:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire T51;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    last = {1{$random}};
    strb = {1{$random}};
    size = {1{$random}};
    data = {2{$random}};
    addr = {1{$random}};
    id = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T4 | T3;
  assign T3 = 3'h3 <= io_aw_bits_size;
  assign T4 = io_aw_valid ^ 1'h1;
  assign io_smi_resp_ready = T5;
  assign T5 = state == 3'h3;
  assign T52 = reset ? 3'h0 : T6;
  assign T6 = T35 ? 3'h0 : T7;
  assign T7 = T34 ? 3'h4 : T8;
  assign T8 = T16 ? T13 : T9;
  assign T9 = T12 ? 3'h2 : T10;
  assign T10 = T11 ? 3'h1 : state;
  assign T11 = io_aw_ready & io_aw_valid;
  assign T12 = io_w_ready & io_w_valid;
  assign T13 = last ? 3'h3 : 3'h1;
  assign T14 = T12 ? io_w_bits_last : T15;
  assign T15 = T11 ? 1'h0 : last;
  assign T16 = T33 & T17;
  assign T17 = strb == 1'h0;
  assign T18 = T28 ? 1'h0 : T19;
  assign T19 = T12 ? T20 : strb;
  assign T20 = T21;
  assign T21 = T22[1'h0:1'h0];
  assign T22 = T23 & T53;
  assign T53 = {248'h0, io_w_bits_strb};
  assign T23 = T24 - 256'h1;
  assign T24 = 1'h1 << T25;
  assign T25 = 1'h1 << size;
  assign T26 = T11 ? io_aw_bits_size : size;
  assign T28 = T33 & T29;
  assign T29 = T32 & T30;
  assign T30 = io_smi_req_ready | T31;
  assign T31 = strb ^ 1'h1;
  assign T32 = T17 ^ 1'h1;
  assign T33 = state == 3'h2;
  assign T34 = io_smi_resp_ready & io_smi_resp_valid;
  assign T35 = io_b_ready & io_b_valid;
  assign io_smi_req_bits_data = data;
  assign T36 = T28 ? 64'h0 : T37;
  assign T37 = T12 ? io_w_bits_data : data;
  assign io_smi_req_bits_addr = addr;
  assign T39 = T28 ? T42 : T40;
  assign T40 = T11 ? T41 : addr;
  assign T41 = io_aw_bits_addr[4'h8:2'h3];
  assign T42 = addr + 6'h1;
  assign io_smi_req_bits_rw = 1'h1;
  assign io_smi_req_valid = T43;
  assign T43 = T44 & strb;
  assign T44 = state == 3'h2;
  assign io_b_bits_user = T45;
  assign T45 = 1'h0;
  assign io_b_bits_id = T46;
  assign T46 = id;
  assign T47 = T11 ? io_aw_bits_id : id;
  assign io_b_bits_resp = T48;
  assign T48 = 2'h0;
  assign io_b_valid = T49;
  assign T49 = state == 3'h4;
  assign io_w_ready = T50;
  assign T50 = state == 3'h1;
  assign io_aw_ready = T51;
  assign T51 = state == 3'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Nasti size must be >= SMI size");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h4;
    end else if(T16) begin
      state <= T13;
    end else if(T12) begin
      state <= 3'h2;
    end else if(T11) begin
      state <= 3'h1;
    end
    if(T12) begin
      last <= io_w_bits_last;
    end else if(T11) begin
      last <= 1'h0;
    end
    if(T28) begin
      strb <= 1'h0;
    end else if(T12) begin
      strb <= T20;
    end
    if(T11) begin
      size <= io_aw_bits_size;
    end
    if(T28) begin
      data <= 64'h0;
    end else if(T12) begin
      data <= io_w_bits_data;
    end
    if(T28) begin
      addr <= T42;
    end else if(T11) begin
      addr <= T41;
    end
    if(T11) begin
      id <= io_aw_bits_id;
    end
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_rw,
    input [5:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_rw,
    input [5:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_rw,
    output[5:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T27;
  wire T3;
  wire T4;
  wire[63:0] T5;
  wire T6;
  wire[5:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T27 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_data = T5;
  assign T5 = T6 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T6 = chosen;
  assign io_out_bits_addr = T7;
  assign T7 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_rw = T8;
  assign T8 = T6 ? io_in_1_bits_rw : io_in_0_bits_rw;
  assign io_out_valid = T9;
  assign T9 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = T18 | T12;
  assign T12 = T13 ^ 1'h1;
  assign T13 = T16 | T14;
  assign T14 = io_in_1_valid & T15;
  assign T15 = last_grant < 1'h1;
  assign T16 = io_in_0_valid & T17;
  assign T17 = last_grant < 1'h0;
  assign T18 = last_grant < 1'h0;
  assign io_in_1_ready = T19;
  assign T19 = T20 & io_out_ready;
  assign T20 = T24 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = T23 | io_in_0_valid;
  assign T23 = T16 | T14;
  assign T24 = T26 & T25;
  assign T25 = last_grant < 1'h1;
  assign T26 = T16 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module SMIArbiter_1(input clk, input reset,
    output io_in_1_req_ready,
    input  io_in_1_req_valid,
    input  io_in_1_req_bits_rw,
    input [5:0] io_in_1_req_bits_addr,
    input [63:0] io_in_1_req_bits_data,
    input  io_in_1_resp_ready,
    output io_in_1_resp_valid,
    output[63:0] io_in_1_resp_bits,
    output io_in_0_req_ready,
    input  io_in_0_req_valid,
    input  io_in_0_req_bits_rw,
    input [5:0] io_in_0_req_bits_addr,
    input [63:0] io_in_0_req_bits_data,
    input  io_in_0_resp_ready,
    output io_in_0_resp_valid,
    output[63:0] io_in_0_resp_bits,
    input  io_out_req_ready,
    output io_out_req_valid,
    output io_out_req_bits_rw,
    output[5:0] io_out_req_bits_addr,
    output[63:0] io_out_req_bits_data,
    output io_out_resp_ready,
    input  io_out_resp_valid,
    input [63:0] io_out_resp_bits
);

  wire T0;
  wire T1;
  reg  wait_resp;
  wire T15;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  choice;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire req_arb_io_in_1_ready;
  wire req_arb_io_in_0_ready;
  wire req_arb_io_out_valid;
  wire req_arb_io_out_bits_rw;
  wire[5:0] req_arb_io_out_bits_addr;
  wire[63:0] req_arb_io_out_bits_data;
  wire req_arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wait_resp = {1{$random}};
    choice = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_out_req_ready & T1;
  assign T1 = wait_resp ^ 1'h1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = T5 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : wait_resp;
  assign T4 = io_out_req_ready & io_out_req_valid;
  assign T5 = io_out_resp_ready & io_out_resp_valid;
  assign io_out_resp_ready = T6;
  assign T6 = T7 ? io_in_1_resp_ready : io_in_0_resp_ready;
  assign T7 = choice;
  assign T8 = T4 ? req_arb_io_chosen : choice;
  assign io_out_req_bits_data = req_arb_io_out_bits_data;
  assign io_out_req_bits_addr = req_arb_io_out_bits_addr;
  assign io_out_req_bits_rw = req_arb_io_out_bits_rw;
  assign io_out_req_valid = T9;
  assign T9 = req_arb_io_out_valid & T10;
  assign T10 = wait_resp ^ 1'h1;
  assign io_in_0_resp_bits = io_out_resp_bits;
  assign io_in_0_resp_valid = T11;
  assign T11 = io_out_resp_valid & T12;
  assign T12 = choice == 1'h0;
  assign io_in_0_req_ready = req_arb_io_in_0_ready;
  assign io_in_1_resp_bits = io_out_resp_bits;
  assign io_in_1_resp_valid = T13;
  assign T13 = io_out_resp_valid & T14;
  assign T14 = choice == 1'h1;
  assign io_in_1_req_ready = req_arb_io_in_1_ready;
  RRArbiter_1 req_arb(.clk(clk), .reset(reset),
       .io_in_1_ready( req_arb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_req_valid ),
       .io_in_1_bits_rw( io_in_1_req_bits_rw ),
       .io_in_1_bits_addr( io_in_1_req_bits_addr ),
       .io_in_1_bits_data( io_in_1_req_bits_data ),
       .io_in_0_ready( req_arb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_req_valid ),
       .io_in_0_bits_rw( io_in_0_req_bits_rw ),
       .io_in_0_bits_addr( io_in_0_req_bits_addr ),
       .io_in_0_bits_data( io_in_0_req_bits_data ),
       .io_out_ready( T0 ),
       .io_out_valid( req_arb_io_out_valid ),
       .io_out_bits_rw( req_arb_io_out_bits_rw ),
       .io_out_bits_addr( req_arb_io_out_bits_addr ),
       .io_out_bits_data( req_arb_io_out_bits_data ),
       .io_chosen( req_arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      wait_resp <= 1'h0;
    end else if(T5) begin
      wait_resp <= 1'h0;
    end else if(T4) begin
      wait_resp <= 1'h1;
    end
    if(T4) begin
      choice <= req_arb_io_chosen;
    end
  end
endmodule

module SMIIONastiIOConverter_1(input clk, input reset,
    output io_nasti_aw_ready,
    input  io_nasti_aw_valid,
    input [31:0] io_nasti_aw_bits_addr,
    input [7:0] io_nasti_aw_bits_len,
    input [2:0] io_nasti_aw_bits_size,
    input [1:0] io_nasti_aw_bits_burst,
    input  io_nasti_aw_bits_lock,
    input [3:0] io_nasti_aw_bits_cache,
    input [2:0] io_nasti_aw_bits_prot,
    input [3:0] io_nasti_aw_bits_qos,
    input [3:0] io_nasti_aw_bits_region,
    input [4:0] io_nasti_aw_bits_id,
    input  io_nasti_aw_bits_user,
    output io_nasti_w_ready,
    input  io_nasti_w_valid,
    input [63:0] io_nasti_w_bits_data,
    input  io_nasti_w_bits_last,
    input [7:0] io_nasti_w_bits_strb,
    input  io_nasti_w_bits_user,
    input  io_nasti_b_ready,
    output io_nasti_b_valid,
    output[1:0] io_nasti_b_bits_resp,
    output[4:0] io_nasti_b_bits_id,
    output io_nasti_b_bits_user,
    output io_nasti_ar_ready,
    input  io_nasti_ar_valid,
    input [31:0] io_nasti_ar_bits_addr,
    input [7:0] io_nasti_ar_bits_len,
    input [2:0] io_nasti_ar_bits_size,
    input [1:0] io_nasti_ar_bits_burst,
    input  io_nasti_ar_bits_lock,
    input [3:0] io_nasti_ar_bits_cache,
    input [2:0] io_nasti_ar_bits_prot,
    input [3:0] io_nasti_ar_bits_qos,
    input [3:0] io_nasti_ar_bits_region,
    input [4:0] io_nasti_ar_bits_id,
    input  io_nasti_ar_bits_user,
    input  io_nasti_r_ready,
    output io_nasti_r_valid,
    output[1:0] io_nasti_r_bits_resp,
    output[63:0] io_nasti_r_bits_data,
    output io_nasti_r_bits_last,
    output[4:0] io_nasti_r_bits_id,
    output io_nasti_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[5:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire reader_io_ar_ready;
  wire reader_io_r_valid;
  wire[1:0] reader_io_r_bits_resp;
  wire[63:0] reader_io_r_bits_data;
  wire reader_io_r_bits_last;
  wire[4:0] reader_io_r_bits_id;
  wire reader_io_r_bits_user;
  wire reader_io_smi_req_valid;
  wire reader_io_smi_req_bits_rw;
  wire[5:0] reader_io_smi_req_bits_addr;
  wire reader_io_smi_resp_ready;
  wire writer_io_aw_ready;
  wire writer_io_w_ready;
  wire writer_io_b_valid;
  wire[1:0] writer_io_b_bits_resp;
  wire[4:0] writer_io_b_bits_id;
  wire writer_io_b_bits_user;
  wire writer_io_smi_req_valid;
  wire writer_io_smi_req_bits_rw;
  wire[5:0] writer_io_smi_req_bits_addr;
  wire[63:0] writer_io_smi_req_bits_data;
  wire writer_io_smi_resp_ready;
  wire arb_io_in_1_req_ready;
  wire arb_io_in_1_resp_valid;
  wire[63:0] arb_io_in_1_resp_bits;
  wire arb_io_in_0_req_ready;
  wire arb_io_in_0_resp_valid;
  wire[63:0] arb_io_in_0_resp_bits;
  wire arb_io_out_req_valid;
  wire arb_io_out_req_bits_rw;
  wire[5:0] arb_io_out_req_bits_addr;
  wire[63:0] arb_io_out_req_bits_data;
  wire arb_io_out_resp_ready;


  assign io_smi_resp_ready = arb_io_out_resp_ready;
  assign io_smi_req_bits_data = arb_io_out_req_bits_data;
  assign io_smi_req_bits_addr = arb_io_out_req_bits_addr;
  assign io_smi_req_bits_rw = arb_io_out_req_bits_rw;
  assign io_smi_req_valid = arb_io_out_req_valid;
  assign io_nasti_r_bits_user = reader_io_r_bits_user;
  assign io_nasti_r_bits_id = reader_io_r_bits_id;
  assign io_nasti_r_bits_last = reader_io_r_bits_last;
  assign io_nasti_r_bits_data = reader_io_r_bits_data;
  assign io_nasti_r_bits_resp = reader_io_r_bits_resp;
  assign io_nasti_r_valid = reader_io_r_valid;
  assign io_nasti_ar_ready = reader_io_ar_ready;
  assign io_nasti_b_bits_user = writer_io_b_bits_user;
  assign io_nasti_b_bits_id = writer_io_b_bits_id;
  assign io_nasti_b_bits_resp = writer_io_b_bits_resp;
  assign io_nasti_b_valid = writer_io_b_valid;
  assign io_nasti_w_ready = writer_io_w_ready;
  assign io_nasti_aw_ready = writer_io_aw_ready;
  SMIIONastiReadIOConverter_1 reader(.clk(clk), .reset(reset),
       .io_ar_ready( reader_io_ar_ready ),
       .io_ar_valid( io_nasti_ar_valid ),
       .io_ar_bits_addr( io_nasti_ar_bits_addr ),
       .io_ar_bits_len( io_nasti_ar_bits_len ),
       .io_ar_bits_size( io_nasti_ar_bits_size ),
       .io_ar_bits_burst( io_nasti_ar_bits_burst ),
       .io_ar_bits_lock( io_nasti_ar_bits_lock ),
       .io_ar_bits_cache( io_nasti_ar_bits_cache ),
       .io_ar_bits_prot( io_nasti_ar_bits_prot ),
       .io_ar_bits_qos( io_nasti_ar_bits_qos ),
       .io_ar_bits_region( io_nasti_ar_bits_region ),
       .io_ar_bits_id( io_nasti_ar_bits_id ),
       .io_ar_bits_user( io_nasti_ar_bits_user ),
       .io_r_ready( io_nasti_r_ready ),
       .io_r_valid( reader_io_r_valid ),
       .io_r_bits_resp( reader_io_r_bits_resp ),
       .io_r_bits_data( reader_io_r_bits_data ),
       .io_r_bits_last( reader_io_r_bits_last ),
       .io_r_bits_id( reader_io_r_bits_id ),
       .io_r_bits_user( reader_io_r_bits_user ),
       .io_smi_req_ready( arb_io_in_0_req_ready ),
       .io_smi_req_valid( reader_io_smi_req_valid ),
       .io_smi_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_smi_req_bits_data(  )
       .io_smi_resp_ready( reader_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_0_resp_valid ),
       .io_smi_resp_bits( arb_io_in_0_resp_bits )
  );
  SMIIONastiWriteIOConverter_1 writer(.clk(clk), .reset(reset),
       .io_aw_ready( writer_io_aw_ready ),
       .io_aw_valid( io_nasti_aw_valid ),
       .io_aw_bits_addr( io_nasti_aw_bits_addr ),
       .io_aw_bits_len( io_nasti_aw_bits_len ),
       .io_aw_bits_size( io_nasti_aw_bits_size ),
       .io_aw_bits_burst( io_nasti_aw_bits_burst ),
       .io_aw_bits_lock( io_nasti_aw_bits_lock ),
       .io_aw_bits_cache( io_nasti_aw_bits_cache ),
       .io_aw_bits_prot( io_nasti_aw_bits_prot ),
       .io_aw_bits_qos( io_nasti_aw_bits_qos ),
       .io_aw_bits_region( io_nasti_aw_bits_region ),
       .io_aw_bits_id( io_nasti_aw_bits_id ),
       .io_aw_bits_user( io_nasti_aw_bits_user ),
       .io_w_ready( writer_io_w_ready ),
       .io_w_valid( io_nasti_w_valid ),
       .io_w_bits_data( io_nasti_w_bits_data ),
       .io_w_bits_last( io_nasti_w_bits_last ),
       .io_w_bits_strb( io_nasti_w_bits_strb ),
       .io_w_bits_user( io_nasti_w_bits_user ),
       .io_b_ready( io_nasti_b_ready ),
       .io_b_valid( writer_io_b_valid ),
       .io_b_bits_resp( writer_io_b_bits_resp ),
       .io_b_bits_id( writer_io_b_bits_id ),
       .io_b_bits_user( writer_io_b_bits_user ),
       .io_smi_req_ready( arb_io_in_1_req_ready ),
       .io_smi_req_valid( writer_io_smi_req_valid ),
       .io_smi_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( writer_io_smi_req_bits_data ),
       .io_smi_resp_ready( writer_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_1_resp_valid ),
       .io_smi_resp_bits( arb_io_in_1_resp_bits )
  );
  SMIArbiter_1 arb(.clk(clk), .reset(reset),
       .io_in_1_req_ready( arb_io_in_1_req_ready ),
       .io_in_1_req_valid( writer_io_smi_req_valid ),
       .io_in_1_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_in_1_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_in_1_req_bits_data( writer_io_smi_req_bits_data ),
       .io_in_1_resp_ready( writer_io_smi_resp_ready ),
       .io_in_1_resp_valid( arb_io_in_1_resp_valid ),
       .io_in_1_resp_bits( arb_io_in_1_resp_bits ),
       .io_in_0_req_ready( arb_io_in_0_req_ready ),
       .io_in_0_req_valid( reader_io_smi_req_valid ),
       .io_in_0_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_in_0_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_in_0_req_bits_data(  )
       .io_in_0_resp_ready( reader_io_smi_resp_ready ),
       .io_in_0_resp_valid( arb_io_in_0_resp_valid ),
       .io_in_0_resp_bits( arb_io_in_0_resp_bits ),
       .io_out_req_ready( io_smi_req_ready ),
       .io_out_req_valid( arb_io_out_req_valid ),
       .io_out_req_bits_rw( arb_io_out_req_bits_rw ),
       .io_out_req_bits_addr( arb_io_out_req_bits_addr ),
       .io_out_req_bits_data( arb_io_out_req_bits_data ),
       .io_out_resp_ready( arb_io_out_resp_ready ),
       .io_out_resp_valid( io_smi_resp_valid ),
       .io_out_resp_bits( io_smi_resp_bits )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign arb.io_in_0_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
endmodule

module OuterMemorySystem(input clk, input reset,
    output io_tiles_cached_0_acquire_ready,
    input  io_tiles_cached_0_acquire_valid,
    input [25:0] io_tiles_cached_0_acquire_bits_addr_block,
    input [1:0] io_tiles_cached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_acquire_bits_addr_beat,
    input  io_tiles_cached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_cached_0_acquire_bits_a_type,
    input [16:0] io_tiles_cached_0_acquire_bits_union,
    input [127:0] io_tiles_cached_0_acquire_bits_data,
    input  io_tiles_cached_0_grant_ready,
    output io_tiles_cached_0_grant_valid,
    output[1:0] io_tiles_cached_0_grant_bits_addr_beat,
    output[1:0] io_tiles_cached_0_grant_bits_client_xact_id,
    output[3:0] io_tiles_cached_0_grant_bits_manager_xact_id,
    output io_tiles_cached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_cached_0_grant_bits_g_type,
    output[127:0] io_tiles_cached_0_grant_bits_data,
    input  io_tiles_cached_0_probe_ready,
    output io_tiles_cached_0_probe_valid,
    output[25:0] io_tiles_cached_0_probe_bits_addr_block,
    output[1:0] io_tiles_cached_0_probe_bits_p_type,
    output io_tiles_cached_0_release_ready,
    input  io_tiles_cached_0_release_valid,
    input [1:0] io_tiles_cached_0_release_bits_addr_beat,
    input [25:0] io_tiles_cached_0_release_bits_addr_block,
    input [1:0] io_tiles_cached_0_release_bits_client_xact_id,
    input [2:0] io_tiles_cached_0_release_bits_r_type,
    input  io_tiles_cached_0_release_bits_voluntary,
    input [127:0] io_tiles_cached_0_release_bits_data,
    output io_tiles_uncached_0_acquire_ready,
    input  io_tiles_uncached_0_acquire_valid,
    input [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
    input [1:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_uncached_0_acquire_bits_addr_beat,
    input  io_tiles_uncached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_uncached_0_acquire_bits_a_type,
    input [16:0] io_tiles_uncached_0_acquire_bits_union,
    input [127:0] io_tiles_uncached_0_acquire_bits_data,
    input  io_tiles_uncached_0_grant_ready,
    output io_tiles_uncached_0_grant_valid,
    output[1:0] io_tiles_uncached_0_grant_bits_addr_beat,
    output[1:0] io_tiles_uncached_0_grant_bits_client_xact_id,
    output[3:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
    output io_tiles_uncached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_uncached_0_grant_bits_g_type,
    output[127:0] io_tiles_uncached_0_grant_bits_data,
    output io_htif_uncached_acquire_ready,
    input  io_htif_uncached_acquire_valid,
    input [25:0] io_htif_uncached_acquire_bits_addr_block,
    input [1:0] io_htif_uncached_acquire_bits_client_xact_id,
    input [1:0] io_htif_uncached_acquire_bits_addr_beat,
    input  io_htif_uncached_acquire_bits_is_builtin_type,
    input [2:0] io_htif_uncached_acquire_bits_a_type,
    input [16:0] io_htif_uncached_acquire_bits_union,
    input [127:0] io_htif_uncached_acquire_bits_data,
    input  io_htif_uncached_grant_ready,
    output io_htif_uncached_grant_valid,
    output[1:0] io_htif_uncached_grant_bits_addr_beat,
    output[1:0] io_htif_uncached_grant_bits_client_xact_id,
    output[3:0] io_htif_uncached_grant_bits_manager_xact_id,
    output io_htif_uncached_grant_bits_is_builtin_type,
    output[3:0] io_htif_uncached_grant_bits_g_type,
    output[127:0] io_htif_uncached_grant_bits_data,
    input  io_incoherent_0,
    input  io_mem_0_aw_ready,
    output io_mem_0_aw_valid,
    output[31:0] io_mem_0_aw_bits_addr,
    output[7:0] io_mem_0_aw_bits_len,
    output[2:0] io_mem_0_aw_bits_size,
    output[1:0] io_mem_0_aw_bits_burst,
    output io_mem_0_aw_bits_lock,
    output[3:0] io_mem_0_aw_bits_cache,
    output[2:0] io_mem_0_aw_bits_prot,
    output[3:0] io_mem_0_aw_bits_qos,
    output[3:0] io_mem_0_aw_bits_region,
    output[4:0] io_mem_0_aw_bits_id,
    output io_mem_0_aw_bits_user,
    input  io_mem_0_w_ready,
    output io_mem_0_w_valid,
    output[63:0] io_mem_0_w_bits_data,
    output io_mem_0_w_bits_last,
    output[7:0] io_mem_0_w_bits_strb,
    output io_mem_0_w_bits_user,
    output io_mem_0_b_ready,
    input  io_mem_0_b_valid,
    input [1:0] io_mem_0_b_bits_resp,
    input [4:0] io_mem_0_b_bits_id,
    input  io_mem_0_b_bits_user,
    input  io_mem_0_ar_ready,
    output io_mem_0_ar_valid,
    output[31:0] io_mem_0_ar_bits_addr,
    output[7:0] io_mem_0_ar_bits_len,
    output[2:0] io_mem_0_ar_bits_size,
    output[1:0] io_mem_0_ar_bits_burst,
    output io_mem_0_ar_bits_lock,
    output[3:0] io_mem_0_ar_bits_cache,
    output[2:0] io_mem_0_ar_bits_prot,
    output[3:0] io_mem_0_ar_bits_qos,
    output[3:0] io_mem_0_ar_bits_region,
    output[4:0] io_mem_0_ar_bits_id,
    output io_mem_0_ar_bits_user,
    output io_mem_0_r_ready,
    input  io_mem_0_r_valid,
    input [1:0] io_mem_0_r_bits_resp,
    input [63:0] io_mem_0_r_bits_data,
    input  io_mem_0_r_bits_last,
    input [4:0] io_mem_0_r_bits_id,
    input  io_mem_0_r_bits_user,
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
    input  io_csr_0_req_ready,
    output io_csr_0_req_valid,
    output io_csr_0_req_bits_rw,
    output[11:0] io_csr_0_req_bits_addr,
    output[63:0] io_csr_0_req_bits_data,
    output io_csr_0_resp_ready,
    input  io_csr_0_resp_valid,
    input [63:0] io_csr_0_resp_bits,
    input  io_scr_req_ready,
    output io_scr_req_valid,
    output io_scr_req_bits_rw,
    output[5:0] io_scr_req_bits_addr,
    output[63:0] io_scr_req_bits_data,
    output io_scr_resp_ready,
    input  io_scr_resp_valid,
    input [63:0] io_scr_resp_bits,
    input  io_mmio_aw_ready,
    output io_mmio_aw_valid,
    output[31:0] io_mmio_aw_bits_addr,
    output[7:0] io_mmio_aw_bits_len,
    output[2:0] io_mmio_aw_bits_size,
    output[1:0] io_mmio_aw_bits_burst,
    output io_mmio_aw_bits_lock,
    output[3:0] io_mmio_aw_bits_cache,
    output[2:0] io_mmio_aw_bits_prot,
    output[3:0] io_mmio_aw_bits_qos,
    output[3:0] io_mmio_aw_bits_region,
    output[4:0] io_mmio_aw_bits_id,
    output io_mmio_aw_bits_user,
    input  io_mmio_w_ready,
    output io_mmio_w_valid,
    output[63:0] io_mmio_w_bits_data,
    output io_mmio_w_bits_last,
    output[7:0] io_mmio_w_bits_strb,
    output io_mmio_w_bits_user,
    output io_mmio_b_ready,
    input  io_mmio_b_valid,
    input [1:0] io_mmio_b_bits_resp,
    input [4:0] io_mmio_b_bits_id,
    input  io_mmio_b_bits_user,
    input  io_mmio_ar_ready,
    output io_mmio_ar_valid,
    output[31:0] io_mmio_ar_bits_addr,
    output[7:0] io_mmio_ar_bits_len,
    output[2:0] io_mmio_ar_bits_size,
    output[1:0] io_mmio_ar_bits_burst,
    output io_mmio_ar_bits_lock,
    output[3:0] io_mmio_ar_bits_cache,
    output[2:0] io_mmio_ar_bits_prot,
    output[3:0] io_mmio_ar_bits_qos,
    output[3:0] io_mmio_ar_bits_region,
    output[4:0] io_mmio_ar_bits_id,
    output io_mmio_ar_bits_user,
    output io_mmio_r_ready,
    input  io_mmio_r_valid,
    input [1:0] io_mmio_r_bits_resp,
    input [63:0] io_mmio_r_bits_data,
    input  io_mmio_r_bits_last,
    input [4:0] io_mmio_r_bits_id,
    input  io_mmio_r_bits_user
);

  wire ClientTileLinkIOWrapper_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOWrapper_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block;
  wire[1:0] ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOWrapper_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_io_out_release_valid;
  wire ClientTileLinkIOWrapper_1_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_1_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_1_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block;
  wire[1:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_1_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_1_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_1_io_out_release_valid;
  wire ClientTileLinkIOWrapper_2_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_2_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat;
  wire[3:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id;
  wire ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_2_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block;
  wire[3:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_2_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_2_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_2_io_out_release_valid;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[31:0] Queue_io_deq_bits_addr;
  wire[7:0] Queue_io_deq_bits_len;
  wire[2:0] Queue_io_deq_bits_size;
  wire[1:0] Queue_io_deq_bits_burst;
  wire Queue_io_deq_bits_lock;
  wire[3:0] Queue_io_deq_bits_cache;
  wire[2:0] Queue_io_deq_bits_prot;
  wire[3:0] Queue_io_deq_bits_qos;
  wire[3:0] Queue_io_deq_bits_region;
  wire[4:0] Queue_io_deq_bits_id;
  wire Queue_io_deq_bits_user;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[31:0] Queue_1_io_deq_bits_addr;
  wire[7:0] Queue_1_io_deq_bits_len;
  wire[2:0] Queue_1_io_deq_bits_size;
  wire[1:0] Queue_1_io_deq_bits_burst;
  wire Queue_1_io_deq_bits_lock;
  wire[3:0] Queue_1_io_deq_bits_cache;
  wire[2:0] Queue_1_io_deq_bits_prot;
  wire[3:0] Queue_1_io_deq_bits_qos;
  wire[3:0] Queue_1_io_deq_bits_region;
  wire[4:0] Queue_1_io_deq_bits_id;
  wire Queue_1_io_deq_bits_user;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire[63:0] Queue_2_io_deq_bits_data;
  wire Queue_2_io_deq_bits_last;
  wire[7:0] Queue_2_io_deq_bits_strb;
  wire Queue_2_io_deq_bits_user;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire[1:0] Queue_3_io_deq_bits_resp;
  wire[63:0] Queue_3_io_deq_bits_data;
  wire Queue_3_io_deq_bits_last;
  wire[4:0] Queue_3_io_deq_bits_id;
  wire Queue_3_io_deq_bits_user;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_resp;
  wire[4:0] Queue_4_io_deq_bits_id;
  wire Queue_4_io_deq_bits_user;
  wire rtc_io_aw_valid;
  wire[31:0] rtc_io_aw_bits_addr;
  wire[7:0] rtc_io_aw_bits_len;
  wire[2:0] rtc_io_aw_bits_size;
  wire[1:0] rtc_io_aw_bits_burst;
  wire rtc_io_aw_bits_lock;
  wire[3:0] rtc_io_aw_bits_cache;
  wire[2:0] rtc_io_aw_bits_prot;
  wire[3:0] rtc_io_aw_bits_qos;
  wire[3:0] rtc_io_aw_bits_region;
  wire[4:0] rtc_io_aw_bits_id;
  wire rtc_io_aw_bits_user;
  wire rtc_io_w_valid;
  wire[63:0] rtc_io_w_bits_data;
  wire rtc_io_w_bits_last;
  wire[7:0] rtc_io_w_bits_strb;
  wire rtc_io_w_bits_user;
  wire rtc_io_b_ready;
  wire rtc_io_ar_valid;
  wire rtc_io_r_ready;
  wire ClientTileLinkIOUnwrapper_io_in_acquire_ready;
  wire ClientTileLinkIOUnwrapper_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_addr_beat;
  wire[3:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_client_xact_id;
  wire ClientTileLinkIOUnwrapper_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOUnwrapper_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_data;
  wire ClientTileLinkIOUnwrapper_io_in_probe_valid;
  wire ClientTileLinkIOUnwrapper_io_in_release_ready;
  wire ClientTileLinkIOUnwrapper_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_block;
  wire[3:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOUnwrapper_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_data;
  wire ClientTileLinkIOUnwrapper_io_out_grant_ready;
  wire TileLinkIONarrower_io_in_acquire_ready;
  wire TileLinkIONarrower_io_in_grant_valid;
  wire[1:0] TileLinkIONarrower_io_in_grant_bits_addr_beat;
  wire[3:0] TileLinkIONarrower_io_in_grant_bits_client_xact_id;
  wire TileLinkIONarrower_io_in_grant_bits_manager_xact_id;
  wire TileLinkIONarrower_io_in_grant_bits_is_builtin_type;
  wire[3:0] TileLinkIONarrower_io_in_grant_bits_g_type;
  wire[127:0] TileLinkIONarrower_io_in_grant_bits_data;
  wire TileLinkIONarrower_io_out_acquire_valid;
  wire[25:0] TileLinkIONarrower_io_out_acquire_bits_addr_block;
  wire[3:0] TileLinkIONarrower_io_out_acquire_bits_client_xact_id;
  wire[2:0] TileLinkIONarrower_io_out_acquire_bits_addr_beat;
  wire TileLinkIONarrower_io_out_acquire_bits_is_builtin_type;
  wire[2:0] TileLinkIONarrower_io_out_acquire_bits_a_type;
  wire[11:0] TileLinkIONarrower_io_out_acquire_bits_union;
  wire[63:0] TileLinkIONarrower_io_out_acquire_bits_data;
  wire TileLinkIONarrower_io_out_grant_ready;
  wire NastiIOTileLinkIOConverter_io_tl_acquire_ready;
  wire NastiIOTileLinkIOConverter_io_tl_grant_valid;
  wire[2:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_addr_beat;
  wire[3:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id;
  wire NastiIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id;
  wire NastiIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type;
  wire[3:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_g_type;
  wire[63:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_data;
  wire NastiIOTileLinkIOConverter_io_nasti_aw_valid;
  wire[31:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_addr;
  wire[7:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_len;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_size;
  wire[1:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_burst;
  wire NastiIOTileLinkIOConverter_io_nasti_aw_bits_lock;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_cache;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_prot;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_qos;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_region;
  wire[4:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_id;
  wire NastiIOTileLinkIOConverter_io_nasti_aw_bits_user;
  wire NastiIOTileLinkIOConverter_io_nasti_w_valid;
  wire[63:0] NastiIOTileLinkIOConverter_io_nasti_w_bits_data;
  wire NastiIOTileLinkIOConverter_io_nasti_w_bits_last;
  wire[7:0] NastiIOTileLinkIOConverter_io_nasti_w_bits_strb;
  wire NastiIOTileLinkIOConverter_io_nasti_w_bits_user;
  wire NastiIOTileLinkIOConverter_io_nasti_b_ready;
  wire NastiIOTileLinkIOConverter_io_nasti_ar_valid;
  wire[31:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_addr;
  wire[7:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_len;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_size;
  wire[1:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_burst;
  wire NastiIOTileLinkIOConverter_io_nasti_ar_bits_lock;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_cache;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_prot;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_qos;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_region;
  wire[4:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_id;
  wire NastiIOTileLinkIOConverter_io_nasti_ar_bits_user;
  wire NastiIOTileLinkIOConverter_io_nasti_r_ready;
  wire L2BroadcastHub_io_inner_acquire_ready;
  wire L2BroadcastHub_io_inner_grant_valid;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_addr_beat;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_client_xact_id;
  wire[3:0] L2BroadcastHub_io_inner_grant_bits_manager_xact_id;
  wire L2BroadcastHub_io_inner_grant_bits_is_builtin_type;
  wire[3:0] L2BroadcastHub_io_inner_grant_bits_g_type;
  wire[127:0] L2BroadcastHub_io_inner_grant_bits_data;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_client_id;
  wire L2BroadcastHub_io_inner_finish_ready;
  wire L2BroadcastHub_io_inner_probe_valid;
  wire[25:0] L2BroadcastHub_io_inner_probe_bits_addr_block;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_p_type;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_client_id;
  wire L2BroadcastHub_io_inner_release_ready;
  wire L2BroadcastHub_io_outer_acquire_valid;
  wire[25:0] L2BroadcastHub_io_outer_acquire_bits_addr_block;
  wire[3:0] L2BroadcastHub_io_outer_acquire_bits_client_xact_id;
  wire[1:0] L2BroadcastHub_io_outer_acquire_bits_addr_beat;
  wire L2BroadcastHub_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] L2BroadcastHub_io_outer_acquire_bits_a_type;
  wire[16:0] L2BroadcastHub_io_outer_acquire_bits_union;
  wire[127:0] L2BroadcastHub_io_outer_acquire_bits_data;
  wire L2BroadcastHub_io_outer_grant_ready;
  wire SMIIONastiIOConverter_io_nasti_aw_ready;
  wire SMIIONastiIOConverter_io_nasti_w_ready;
  wire SMIIONastiIOConverter_io_nasti_b_valid;
  wire[1:0] SMIIONastiIOConverter_io_nasti_b_bits_resp;
  wire[4:0] SMIIONastiIOConverter_io_nasti_b_bits_id;
  wire SMIIONastiIOConverter_io_nasti_b_bits_user;
  wire SMIIONastiIOConverter_io_nasti_ar_ready;
  wire SMIIONastiIOConverter_io_nasti_r_valid;
  wire[1:0] SMIIONastiIOConverter_io_nasti_r_bits_resp;
  wire[63:0] SMIIONastiIOConverter_io_nasti_r_bits_data;
  wire SMIIONastiIOConverter_io_nasti_r_bits_last;
  wire[4:0] SMIIONastiIOConverter_io_nasti_r_bits_id;
  wire SMIIONastiIOConverter_io_nasti_r_bits_user;
  wire SMIIONastiIOConverter_io_smi_req_valid;
  wire SMIIONastiIOConverter_io_smi_req_bits_rw;
  wire[11:0] SMIIONastiIOConverter_io_smi_req_bits_addr;
  wire[63:0] SMIIONastiIOConverter_io_smi_req_bits_data;
  wire SMIIONastiIOConverter_io_smi_resp_ready;
  wire conv_io_nasti_aw_ready;
  wire conv_io_nasti_w_ready;
  wire conv_io_nasti_b_valid;
  wire[1:0] conv_io_nasti_b_bits_resp;
  wire[4:0] conv_io_nasti_b_bits_id;
  wire conv_io_nasti_b_bits_user;
  wire conv_io_nasti_ar_ready;
  wire conv_io_nasti_r_valid;
  wire[1:0] conv_io_nasti_r_bits_resp;
  wire[63:0] conv_io_nasti_r_bits_data;
  wire conv_io_nasti_r_bits_last;
  wire[4:0] conv_io_nasti_r_bits_id;
  wire conv_io_nasti_r_bits_user;
  wire conv_io_smi_req_valid;
  wire conv_io_smi_req_bits_rw;
  wire[5:0] conv_io_smi_req_bits_addr;
  wire[63:0] conv_io_smi_req_bits_data;
  wire conv_io_smi_resp_ready;
  wire l1tol2net_io_clients_2_acquire_ready;
  wire l1tol2net_io_clients_2_grant_valid;
  wire[1:0] l1tol2net_io_clients_2_grant_bits_addr_beat;
  wire[1:0] l1tol2net_io_clients_2_grant_bits_client_xact_id;
  wire[3:0] l1tol2net_io_clients_2_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_2_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_2_grant_bits_g_type;
  wire[127:0] l1tol2net_io_clients_2_grant_bits_data;
  wire l1tol2net_io_clients_2_probe_valid;
  wire[25:0] l1tol2net_io_clients_2_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_2_probe_bits_p_type;
  wire l1tol2net_io_clients_2_release_ready;
  wire l1tol2net_io_clients_1_acquire_ready;
  wire l1tol2net_io_clients_1_grant_valid;
  wire[1:0] l1tol2net_io_clients_1_grant_bits_addr_beat;
  wire[1:0] l1tol2net_io_clients_1_grant_bits_client_xact_id;
  wire[3:0] l1tol2net_io_clients_1_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_1_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_1_grant_bits_g_type;
  wire[127:0] l1tol2net_io_clients_1_grant_bits_data;
  wire l1tol2net_io_clients_1_probe_valid;
  wire[25:0] l1tol2net_io_clients_1_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_1_probe_bits_p_type;
  wire l1tol2net_io_clients_1_release_ready;
  wire l1tol2net_io_clients_0_acquire_ready;
  wire l1tol2net_io_clients_0_grant_valid;
  wire[1:0] l1tol2net_io_clients_0_grant_bits_addr_beat;
  wire[1:0] l1tol2net_io_clients_0_grant_bits_client_xact_id;
  wire[3:0] l1tol2net_io_clients_0_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_0_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_0_grant_bits_g_type;
  wire[127:0] l1tol2net_io_clients_0_grant_bits_data;
  wire l1tol2net_io_clients_0_probe_valid;
  wire[25:0] l1tol2net_io_clients_0_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_0_probe_bits_p_type;
  wire l1tol2net_io_clients_0_release_ready;
  wire l1tol2net_io_managers_0_acquire_valid;
  wire[25:0] l1tol2net_io_managers_0_acquire_bits_addr_block;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_addr_beat;
  wire l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  wire[2:0] l1tol2net_io_managers_0_acquire_bits_a_type;
  wire[16:0] l1tol2net_io_managers_0_acquire_bits_union;
  wire[127:0] l1tol2net_io_managers_0_acquire_bits_data;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_client_id;
  wire l1tol2net_io_managers_0_grant_ready;
  wire l1tol2net_io_managers_0_finish_valid;
  wire[3:0] l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  wire l1tol2net_io_managers_0_probe_ready;
  wire l1tol2net_io_managers_0_release_valid;
  wire[1:0] l1tol2net_io_managers_0_release_bits_addr_beat;
  wire[25:0] l1tol2net_io_managers_0_release_bits_addr_block;
  wire[1:0] l1tol2net_io_managers_0_release_bits_client_xact_id;
  wire[2:0] l1tol2net_io_managers_0_release_bits_r_type;
  wire l1tol2net_io_managers_0_release_bits_voluntary;
  wire[127:0] l1tol2net_io_managers_0_release_bits_data;
  wire[1:0] l1tol2net_io_managers_0_release_bits_client_id;
  wire interconnect_io_masters_1_aw_ready;
  wire interconnect_io_masters_1_w_ready;
  wire interconnect_io_masters_1_b_valid;
  wire[1:0] interconnect_io_masters_1_b_bits_resp;
  wire[4:0] interconnect_io_masters_1_b_bits_id;
  wire interconnect_io_masters_1_b_bits_user;
  wire interconnect_io_masters_1_ar_ready;
  wire interconnect_io_masters_1_r_valid;
  wire[1:0] interconnect_io_masters_1_r_bits_resp;
  wire[63:0] interconnect_io_masters_1_r_bits_data;
  wire interconnect_io_masters_1_r_bits_last;
  wire[4:0] interconnect_io_masters_1_r_bits_id;
  wire interconnect_io_masters_1_r_bits_user;
  wire interconnect_io_masters_0_aw_ready;
  wire interconnect_io_masters_0_w_ready;
  wire interconnect_io_masters_0_b_valid;
  wire[1:0] interconnect_io_masters_0_b_bits_resp;
  wire[4:0] interconnect_io_masters_0_b_bits_id;
  wire interconnect_io_masters_0_b_bits_user;
  wire interconnect_io_masters_0_ar_ready;
  wire interconnect_io_masters_0_r_valid;
  wire[1:0] interconnect_io_masters_0_r_bits_resp;
  wire[63:0] interconnect_io_masters_0_r_bits_data;
  wire interconnect_io_masters_0_r_bits_last;
  wire[4:0] interconnect_io_masters_0_r_bits_id;
  wire interconnect_io_masters_0_r_bits_user;
  wire interconnect_io_slaves_3_aw_valid;
  wire[31:0] interconnect_io_slaves_3_aw_bits_addr;
  wire[7:0] interconnect_io_slaves_3_aw_bits_len;
  wire[2:0] interconnect_io_slaves_3_aw_bits_size;
  wire[1:0] interconnect_io_slaves_3_aw_bits_burst;
  wire interconnect_io_slaves_3_aw_bits_lock;
  wire[3:0] interconnect_io_slaves_3_aw_bits_cache;
  wire[2:0] interconnect_io_slaves_3_aw_bits_prot;
  wire[3:0] interconnect_io_slaves_3_aw_bits_qos;
  wire[3:0] interconnect_io_slaves_3_aw_bits_region;
  wire[4:0] interconnect_io_slaves_3_aw_bits_id;
  wire interconnect_io_slaves_3_aw_bits_user;
  wire interconnect_io_slaves_3_w_valid;
  wire[63:0] interconnect_io_slaves_3_w_bits_data;
  wire interconnect_io_slaves_3_w_bits_last;
  wire[7:0] interconnect_io_slaves_3_w_bits_strb;
  wire interconnect_io_slaves_3_w_bits_user;
  wire interconnect_io_slaves_3_b_ready;
  wire interconnect_io_slaves_3_ar_valid;
  wire[31:0] interconnect_io_slaves_3_ar_bits_addr;
  wire[7:0] interconnect_io_slaves_3_ar_bits_len;
  wire[2:0] interconnect_io_slaves_3_ar_bits_size;
  wire[1:0] interconnect_io_slaves_3_ar_bits_burst;
  wire interconnect_io_slaves_3_ar_bits_lock;
  wire[3:0] interconnect_io_slaves_3_ar_bits_cache;
  wire[2:0] interconnect_io_slaves_3_ar_bits_prot;
  wire[3:0] interconnect_io_slaves_3_ar_bits_qos;
  wire[3:0] interconnect_io_slaves_3_ar_bits_region;
  wire[4:0] interconnect_io_slaves_3_ar_bits_id;
  wire interconnect_io_slaves_3_ar_bits_user;
  wire interconnect_io_slaves_3_r_ready;
  wire interconnect_io_slaves_2_aw_valid;
  wire[31:0] interconnect_io_slaves_2_aw_bits_addr;
  wire[7:0] interconnect_io_slaves_2_aw_bits_len;
  wire[2:0] interconnect_io_slaves_2_aw_bits_size;
  wire[1:0] interconnect_io_slaves_2_aw_bits_burst;
  wire interconnect_io_slaves_2_aw_bits_lock;
  wire[3:0] interconnect_io_slaves_2_aw_bits_cache;
  wire[2:0] interconnect_io_slaves_2_aw_bits_prot;
  wire[3:0] interconnect_io_slaves_2_aw_bits_qos;
  wire[3:0] interconnect_io_slaves_2_aw_bits_region;
  wire[4:0] interconnect_io_slaves_2_aw_bits_id;
  wire interconnect_io_slaves_2_aw_bits_user;
  wire interconnect_io_slaves_2_w_valid;
  wire[63:0] interconnect_io_slaves_2_w_bits_data;
  wire interconnect_io_slaves_2_w_bits_last;
  wire[7:0] interconnect_io_slaves_2_w_bits_strb;
  wire interconnect_io_slaves_2_w_bits_user;
  wire interconnect_io_slaves_2_b_ready;
  wire interconnect_io_slaves_2_ar_valid;
  wire[31:0] interconnect_io_slaves_2_ar_bits_addr;
  wire[7:0] interconnect_io_slaves_2_ar_bits_len;
  wire[2:0] interconnect_io_slaves_2_ar_bits_size;
  wire[1:0] interconnect_io_slaves_2_ar_bits_burst;
  wire interconnect_io_slaves_2_ar_bits_lock;
  wire[3:0] interconnect_io_slaves_2_ar_bits_cache;
  wire[2:0] interconnect_io_slaves_2_ar_bits_prot;
  wire[3:0] interconnect_io_slaves_2_ar_bits_qos;
  wire[3:0] interconnect_io_slaves_2_ar_bits_region;
  wire[4:0] interconnect_io_slaves_2_ar_bits_id;
  wire interconnect_io_slaves_2_ar_bits_user;
  wire interconnect_io_slaves_2_r_ready;
  wire interconnect_io_slaves_1_aw_valid;
  wire[31:0] interconnect_io_slaves_1_aw_bits_addr;
  wire[7:0] interconnect_io_slaves_1_aw_bits_len;
  wire[2:0] interconnect_io_slaves_1_aw_bits_size;
  wire[1:0] interconnect_io_slaves_1_aw_bits_burst;
  wire interconnect_io_slaves_1_aw_bits_lock;
  wire[3:0] interconnect_io_slaves_1_aw_bits_cache;
  wire[2:0] interconnect_io_slaves_1_aw_bits_prot;
  wire[3:0] interconnect_io_slaves_1_aw_bits_qos;
  wire[3:0] interconnect_io_slaves_1_aw_bits_region;
  wire[4:0] interconnect_io_slaves_1_aw_bits_id;
  wire interconnect_io_slaves_1_aw_bits_user;
  wire interconnect_io_slaves_1_w_valid;
  wire[63:0] interconnect_io_slaves_1_w_bits_data;
  wire interconnect_io_slaves_1_w_bits_last;
  wire[7:0] interconnect_io_slaves_1_w_bits_strb;
  wire interconnect_io_slaves_1_w_bits_user;
  wire interconnect_io_slaves_1_b_ready;
  wire interconnect_io_slaves_1_ar_valid;
  wire[31:0] interconnect_io_slaves_1_ar_bits_addr;
  wire[7:0] interconnect_io_slaves_1_ar_bits_len;
  wire[2:0] interconnect_io_slaves_1_ar_bits_size;
  wire[1:0] interconnect_io_slaves_1_ar_bits_burst;
  wire interconnect_io_slaves_1_ar_bits_lock;
  wire[3:0] interconnect_io_slaves_1_ar_bits_cache;
  wire[2:0] interconnect_io_slaves_1_ar_bits_prot;
  wire[3:0] interconnect_io_slaves_1_ar_bits_qos;
  wire[3:0] interconnect_io_slaves_1_ar_bits_region;
  wire[4:0] interconnect_io_slaves_1_ar_bits_id;
  wire interconnect_io_slaves_1_ar_bits_user;
  wire interconnect_io_slaves_1_r_ready;
  wire interconnect_io_slaves_0_aw_valid;
  wire[31:0] interconnect_io_slaves_0_aw_bits_addr;
  wire[7:0] interconnect_io_slaves_0_aw_bits_len;
  wire[2:0] interconnect_io_slaves_0_aw_bits_size;
  wire[1:0] interconnect_io_slaves_0_aw_bits_burst;
  wire interconnect_io_slaves_0_aw_bits_lock;
  wire[3:0] interconnect_io_slaves_0_aw_bits_cache;
  wire[2:0] interconnect_io_slaves_0_aw_bits_prot;
  wire[3:0] interconnect_io_slaves_0_aw_bits_qos;
  wire[3:0] interconnect_io_slaves_0_aw_bits_region;
  wire[4:0] interconnect_io_slaves_0_aw_bits_id;
  wire interconnect_io_slaves_0_aw_bits_user;
  wire interconnect_io_slaves_0_w_valid;
  wire[63:0] interconnect_io_slaves_0_w_bits_data;
  wire interconnect_io_slaves_0_w_bits_last;
  wire[7:0] interconnect_io_slaves_0_w_bits_strb;
  wire interconnect_io_slaves_0_w_bits_user;
  wire interconnect_io_slaves_0_b_ready;
  wire interconnect_io_slaves_0_ar_valid;
  wire[31:0] interconnect_io_slaves_0_ar_bits_addr;
  wire[7:0] interconnect_io_slaves_0_ar_bits_len;
  wire[2:0] interconnect_io_slaves_0_ar_bits_size;
  wire[1:0] interconnect_io_slaves_0_ar_bits_burst;
  wire interconnect_io_slaves_0_ar_bits_lock;
  wire[3:0] interconnect_io_slaves_0_ar_bits_cache;
  wire[2:0] interconnect_io_slaves_0_ar_bits_prot;
  wire[3:0] interconnect_io_slaves_0_ar_bits_qos;
  wire[3:0] interconnect_io_slaves_0_ar_bits_region;
  wire[4:0] interconnect_io_slaves_0_ar_bits_id;
  wire interconnect_io_slaves_0_ar_bits_user;
  wire interconnect_io_slaves_0_r_ready;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_backup_req_bits = {1{$random}};
//  assign io_mem_backup_req_valid = {1{$random}};
// synthesis translate_on
`endif
  assign io_mmio_r_ready = interconnect_io_slaves_3_r_ready;
  assign io_mmio_ar_bits_user = interconnect_io_slaves_3_ar_bits_user;
  assign io_mmio_ar_bits_id = interconnect_io_slaves_3_ar_bits_id;
  assign io_mmio_ar_bits_region = interconnect_io_slaves_3_ar_bits_region;
  assign io_mmio_ar_bits_qos = interconnect_io_slaves_3_ar_bits_qos;
  assign io_mmio_ar_bits_prot = interconnect_io_slaves_3_ar_bits_prot;
  assign io_mmio_ar_bits_cache = interconnect_io_slaves_3_ar_bits_cache;
  assign io_mmio_ar_bits_lock = interconnect_io_slaves_3_ar_bits_lock;
  assign io_mmio_ar_bits_burst = interconnect_io_slaves_3_ar_bits_burst;
  assign io_mmio_ar_bits_size = interconnect_io_slaves_3_ar_bits_size;
  assign io_mmio_ar_bits_len = interconnect_io_slaves_3_ar_bits_len;
  assign io_mmio_ar_bits_addr = interconnect_io_slaves_3_ar_bits_addr;
  assign io_mmio_ar_valid = interconnect_io_slaves_3_ar_valid;
  assign io_mmio_b_ready = interconnect_io_slaves_3_b_ready;
  assign io_mmio_w_bits_user = interconnect_io_slaves_3_w_bits_user;
  assign io_mmio_w_bits_strb = interconnect_io_slaves_3_w_bits_strb;
  assign io_mmio_w_bits_last = interconnect_io_slaves_3_w_bits_last;
  assign io_mmio_w_bits_data = interconnect_io_slaves_3_w_bits_data;
  assign io_mmio_w_valid = interconnect_io_slaves_3_w_valid;
  assign io_mmio_aw_bits_user = interconnect_io_slaves_3_aw_bits_user;
  assign io_mmio_aw_bits_id = interconnect_io_slaves_3_aw_bits_id;
  assign io_mmio_aw_bits_region = interconnect_io_slaves_3_aw_bits_region;
  assign io_mmio_aw_bits_qos = interconnect_io_slaves_3_aw_bits_qos;
  assign io_mmio_aw_bits_prot = interconnect_io_slaves_3_aw_bits_prot;
  assign io_mmio_aw_bits_cache = interconnect_io_slaves_3_aw_bits_cache;
  assign io_mmio_aw_bits_lock = interconnect_io_slaves_3_aw_bits_lock;
  assign io_mmio_aw_bits_burst = interconnect_io_slaves_3_aw_bits_burst;
  assign io_mmio_aw_bits_size = interconnect_io_slaves_3_aw_bits_size;
  assign io_mmio_aw_bits_len = interconnect_io_slaves_3_aw_bits_len;
  assign io_mmio_aw_bits_addr = interconnect_io_slaves_3_aw_bits_addr;
  assign io_mmio_aw_valid = interconnect_io_slaves_3_aw_valid;
  assign io_scr_resp_ready = conv_io_smi_resp_ready;
  assign io_scr_req_bits_data = conv_io_smi_req_bits_data;
  assign io_scr_req_bits_addr = conv_io_smi_req_bits_addr;
  assign io_scr_req_bits_rw = conv_io_smi_req_bits_rw;
  assign io_scr_req_valid = conv_io_smi_req_valid;
  assign io_csr_0_resp_ready = SMIIONastiIOConverter_io_smi_resp_ready;
  assign io_csr_0_req_bits_data = SMIIONastiIOConverter_io_smi_req_bits_data;
  assign io_csr_0_req_bits_addr = SMIIONastiIOConverter_io_smi_req_bits_addr;
  assign io_csr_0_req_bits_rw = SMIIONastiIOConverter_io_smi_req_bits_rw;
  assign io_csr_0_req_valid = SMIIONastiIOConverter_io_smi_req_valid;
  assign io_mem_0_r_ready = interconnect_io_slaves_0_r_ready;
  assign io_mem_0_ar_bits_user = interconnect_io_slaves_0_ar_bits_user;
  assign io_mem_0_ar_bits_id = interconnect_io_slaves_0_ar_bits_id;
  assign io_mem_0_ar_bits_region = interconnect_io_slaves_0_ar_bits_region;
  assign io_mem_0_ar_bits_qos = interconnect_io_slaves_0_ar_bits_qos;
  assign io_mem_0_ar_bits_prot = interconnect_io_slaves_0_ar_bits_prot;
  assign io_mem_0_ar_bits_cache = interconnect_io_slaves_0_ar_bits_cache;
  assign io_mem_0_ar_bits_lock = interconnect_io_slaves_0_ar_bits_lock;
  assign io_mem_0_ar_bits_burst = interconnect_io_slaves_0_ar_bits_burst;
  assign io_mem_0_ar_bits_size = interconnect_io_slaves_0_ar_bits_size;
  assign io_mem_0_ar_bits_len = interconnect_io_slaves_0_ar_bits_len;
  assign io_mem_0_ar_bits_addr = interconnect_io_slaves_0_ar_bits_addr;
  assign io_mem_0_ar_valid = interconnect_io_slaves_0_ar_valid;
  assign io_mem_0_b_ready = interconnect_io_slaves_0_b_ready;
  assign io_mem_0_w_bits_user = interconnect_io_slaves_0_w_bits_user;
  assign io_mem_0_w_bits_strb = interconnect_io_slaves_0_w_bits_strb;
  assign io_mem_0_w_bits_last = interconnect_io_slaves_0_w_bits_last;
  assign io_mem_0_w_bits_data = interconnect_io_slaves_0_w_bits_data;
  assign io_mem_0_w_valid = interconnect_io_slaves_0_w_valid;
  assign io_mem_0_aw_bits_user = interconnect_io_slaves_0_aw_bits_user;
  assign io_mem_0_aw_bits_id = interconnect_io_slaves_0_aw_bits_id;
  assign io_mem_0_aw_bits_region = interconnect_io_slaves_0_aw_bits_region;
  assign io_mem_0_aw_bits_qos = interconnect_io_slaves_0_aw_bits_qos;
  assign io_mem_0_aw_bits_prot = interconnect_io_slaves_0_aw_bits_prot;
  assign io_mem_0_aw_bits_cache = interconnect_io_slaves_0_aw_bits_cache;
  assign io_mem_0_aw_bits_lock = interconnect_io_slaves_0_aw_bits_lock;
  assign io_mem_0_aw_bits_burst = interconnect_io_slaves_0_aw_bits_burst;
  assign io_mem_0_aw_bits_size = interconnect_io_slaves_0_aw_bits_size;
  assign io_mem_0_aw_bits_len = interconnect_io_slaves_0_aw_bits_len;
  assign io_mem_0_aw_bits_addr = interconnect_io_slaves_0_aw_bits_addr;
  assign io_mem_0_aw_valid = interconnect_io_slaves_0_aw_valid;
  assign io_htif_uncached_grant_bits_data = ClientTileLinkIOWrapper_1_io_in_grant_bits_data;
  assign io_htif_uncached_grant_bits_g_type = ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type;
  assign io_htif_uncached_grant_bits_is_builtin_type = ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type;
  assign io_htif_uncached_grant_bits_manager_xact_id = ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id;
  assign io_htif_uncached_grant_bits_client_xact_id = ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id;
  assign io_htif_uncached_grant_bits_addr_beat = ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat;
  assign io_htif_uncached_grant_valid = ClientTileLinkIOWrapper_1_io_in_grant_valid;
  assign io_htif_uncached_acquire_ready = ClientTileLinkIOWrapper_1_io_in_acquire_ready;
  assign io_tiles_uncached_0_grant_bits_data = ClientTileLinkIOWrapper_io_in_grant_bits_data;
  assign io_tiles_uncached_0_grant_bits_g_type = ClientTileLinkIOWrapper_io_in_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_addr_beat = ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_valid = ClientTileLinkIOWrapper_io_in_grant_valid;
  assign io_tiles_uncached_0_acquire_ready = ClientTileLinkIOWrapper_io_in_acquire_ready;
  assign io_tiles_cached_0_release_ready = l1tol2net_io_clients_0_release_ready;
  assign io_tiles_cached_0_probe_bits_p_type = l1tol2net_io_clients_0_probe_bits_p_type;
  assign io_tiles_cached_0_probe_bits_addr_block = l1tol2net_io_clients_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_valid = l1tol2net_io_clients_0_probe_valid;
  assign io_tiles_cached_0_grant_bits_data = l1tol2net_io_clients_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_g_type = l1tol2net_io_clients_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_client_xact_id = l1tol2net_io_clients_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_addr_beat = l1tol2net_io_clients_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_valid = l1tol2net_io_clients_0_grant_valid;
  assign io_tiles_cached_0_acquire_ready = l1tol2net_io_clients_0_acquire_ready;
  ClientTileLinkIOWrapper_0 ClientTileLinkIOWrapper(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_io_in_acquire_ready ),
       .io_in_acquire_valid( io_tiles_uncached_0_acquire_valid ),
       .io_in_acquire_bits_addr_block( io_tiles_uncached_0_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( io_tiles_uncached_0_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( io_tiles_uncached_0_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( io_tiles_uncached_0_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( io_tiles_uncached_0_acquire_bits_a_type ),
       .io_in_acquire_bits_union( io_tiles_uncached_0_acquire_bits_union ),
       .io_in_acquire_bits_data( io_tiles_uncached_0_acquire_bits_data ),
       .io_in_grant_ready( io_tiles_uncached_0_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_io_in_grant_bits_data ),
       .io_out_acquire_ready( l1tol2net_io_clients_1_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_io_out_grant_ready ),
       .io_out_grant_valid( l1tol2net_io_clients_1_grant_valid ),
       .io_out_grant_bits_addr_beat( l1tol2net_io_clients_1_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( l1tol2net_io_clients_1_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( l1tol2net_io_clients_1_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( l1tol2net_io_clients_1_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( l1tol2net_io_clients_1_grant_bits_g_type ),
       .io_out_grant_bits_data( l1tol2net_io_clients_1_grant_bits_data ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_io_out_probe_ready ),
       .io_out_probe_valid( l1tol2net_io_clients_1_probe_valid ),
       .io_out_probe_bits_addr_block( l1tol2net_io_clients_1_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( l1tol2net_io_clients_1_probe_bits_p_type ),
       .io_out_release_ready( l1tol2net_io_clients_1_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_io_out_release_valid )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_data(  )
  );
  ClientTileLinkIOWrapper_0 ClientTileLinkIOWrapper_1(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_1_io_in_acquire_ready ),
       .io_in_acquire_valid( io_htif_uncached_acquire_valid ),
       .io_in_acquire_bits_addr_block( io_htif_uncached_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( io_htif_uncached_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( io_htif_uncached_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( io_htif_uncached_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( io_htif_uncached_acquire_bits_a_type ),
       .io_in_acquire_bits_union( io_htif_uncached_acquire_bits_union ),
       .io_in_acquire_bits_data( io_htif_uncached_acquire_bits_data ),
       .io_in_grant_ready( io_htif_uncached_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_1_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_1_io_in_grant_bits_data ),
       .io_out_acquire_ready( l1tol2net_io_clients_2_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_1_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_1_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_1_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_1_io_out_grant_ready ),
       .io_out_grant_valid( l1tol2net_io_clients_2_grant_valid ),
       .io_out_grant_bits_addr_beat( l1tol2net_io_clients_2_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( l1tol2net_io_clients_2_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( l1tol2net_io_clients_2_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( l1tol2net_io_clients_2_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( l1tol2net_io_clients_2_grant_bits_g_type ),
       .io_out_grant_bits_data( l1tol2net_io_clients_2_grant_bits_data ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_1_io_out_probe_ready ),
       .io_out_probe_valid( l1tol2net_io_clients_2_probe_valid ),
       .io_out_probe_bits_addr_block( l1tol2net_io_clients_2_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( l1tol2net_io_clients_2_probe_bits_p_type ),
       .io_out_release_ready( l1tol2net_io_clients_2_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_1_io_out_release_valid )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_data(  )
  );
  RocketChipTileLinkArbiter l1tol2net(.clk(clk), .reset(reset),
       .io_clients_2_acquire_ready( l1tol2net_io_clients_2_acquire_ready ),
       .io_clients_2_acquire_valid( ClientTileLinkIOWrapper_1_io_out_acquire_valid ),
       .io_clients_2_acquire_bits_addr_block( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block ),
       .io_clients_2_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id ),
       .io_clients_2_acquire_bits_addr_beat( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat ),
       .io_clients_2_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type ),
       .io_clients_2_acquire_bits_a_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type ),
       .io_clients_2_acquire_bits_union( ClientTileLinkIOWrapper_1_io_out_acquire_bits_union ),
       .io_clients_2_acquire_bits_data( ClientTileLinkIOWrapper_1_io_out_acquire_bits_data ),
       .io_clients_2_grant_ready( ClientTileLinkIOWrapper_1_io_out_grant_ready ),
       .io_clients_2_grant_valid( l1tol2net_io_clients_2_grant_valid ),
       .io_clients_2_grant_bits_addr_beat( l1tol2net_io_clients_2_grant_bits_addr_beat ),
       .io_clients_2_grant_bits_client_xact_id( l1tol2net_io_clients_2_grant_bits_client_xact_id ),
       .io_clients_2_grant_bits_manager_xact_id( l1tol2net_io_clients_2_grant_bits_manager_xact_id ),
       .io_clients_2_grant_bits_is_builtin_type( l1tol2net_io_clients_2_grant_bits_is_builtin_type ),
       .io_clients_2_grant_bits_g_type( l1tol2net_io_clients_2_grant_bits_g_type ),
       .io_clients_2_grant_bits_data( l1tol2net_io_clients_2_grant_bits_data ),
       .io_clients_2_probe_ready( ClientTileLinkIOWrapper_1_io_out_probe_ready ),
       .io_clients_2_probe_valid( l1tol2net_io_clients_2_probe_valid ),
       .io_clients_2_probe_bits_addr_block( l1tol2net_io_clients_2_probe_bits_addr_block ),
       .io_clients_2_probe_bits_p_type( l1tol2net_io_clients_2_probe_bits_p_type ),
       .io_clients_2_release_ready( l1tol2net_io_clients_2_release_ready ),
       .io_clients_2_release_valid( ClientTileLinkIOWrapper_1_io_out_release_valid ),
       //.io_clients_2_release_bits_addr_beat(  )
       //.io_clients_2_release_bits_addr_block(  )
       //.io_clients_2_release_bits_client_xact_id(  )
       //.io_clients_2_release_bits_r_type(  )
       //.io_clients_2_release_bits_voluntary(  )
       //.io_clients_2_release_bits_data(  )
       .io_clients_1_acquire_ready( l1tol2net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( ClientTileLinkIOWrapper_io_out_acquire_valid ),
       .io_clients_1_acquire_bits_addr_block( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block ),
       .io_clients_1_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id ),
       .io_clients_1_acquire_bits_addr_beat( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat ),
       .io_clients_1_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type ),
       .io_clients_1_acquire_bits_a_type( ClientTileLinkIOWrapper_io_out_acquire_bits_a_type ),
       .io_clients_1_acquire_bits_union( ClientTileLinkIOWrapper_io_out_acquire_bits_union ),
       .io_clients_1_acquire_bits_data( ClientTileLinkIOWrapper_io_out_acquire_bits_data ),
       .io_clients_1_grant_ready( ClientTileLinkIOWrapper_io_out_grant_ready ),
       .io_clients_1_grant_valid( l1tol2net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_addr_beat( l1tol2net_io_clients_1_grant_bits_addr_beat ),
       .io_clients_1_grant_bits_client_xact_id( l1tol2net_io_clients_1_grant_bits_client_xact_id ),
       .io_clients_1_grant_bits_manager_xact_id( l1tol2net_io_clients_1_grant_bits_manager_xact_id ),
       .io_clients_1_grant_bits_is_builtin_type( l1tol2net_io_clients_1_grant_bits_is_builtin_type ),
       .io_clients_1_grant_bits_g_type( l1tol2net_io_clients_1_grant_bits_g_type ),
       .io_clients_1_grant_bits_data( l1tol2net_io_clients_1_grant_bits_data ),
       .io_clients_1_probe_ready( ClientTileLinkIOWrapper_io_out_probe_ready ),
       .io_clients_1_probe_valid( l1tol2net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_addr_block( l1tol2net_io_clients_1_probe_bits_addr_block ),
       .io_clients_1_probe_bits_p_type( l1tol2net_io_clients_1_probe_bits_p_type ),
       .io_clients_1_release_ready( l1tol2net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( ClientTileLinkIOWrapper_io_out_release_valid ),
       //.io_clients_1_release_bits_addr_beat(  )
       //.io_clients_1_release_bits_addr_block(  )
       //.io_clients_1_release_bits_client_xact_id(  )
       //.io_clients_1_release_bits_r_type(  )
       //.io_clients_1_release_bits_voluntary(  )
       //.io_clients_1_release_bits_data(  )
       .io_clients_0_acquire_ready( l1tol2net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_cached_0_acquire_valid ),
       .io_clients_0_acquire_bits_addr_block( io_tiles_cached_0_acquire_bits_addr_block ),
       .io_clients_0_acquire_bits_client_xact_id( io_tiles_cached_0_acquire_bits_client_xact_id ),
       .io_clients_0_acquire_bits_addr_beat( io_tiles_cached_0_acquire_bits_addr_beat ),
       .io_clients_0_acquire_bits_is_builtin_type( io_tiles_cached_0_acquire_bits_is_builtin_type ),
       .io_clients_0_acquire_bits_a_type( io_tiles_cached_0_acquire_bits_a_type ),
       .io_clients_0_acquire_bits_union( io_tiles_cached_0_acquire_bits_union ),
       .io_clients_0_acquire_bits_data( io_tiles_cached_0_acquire_bits_data ),
       .io_clients_0_grant_ready( io_tiles_cached_0_grant_ready ),
       .io_clients_0_grant_valid( l1tol2net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_addr_beat( l1tol2net_io_clients_0_grant_bits_addr_beat ),
       .io_clients_0_grant_bits_client_xact_id( l1tol2net_io_clients_0_grant_bits_client_xact_id ),
       .io_clients_0_grant_bits_manager_xact_id( l1tol2net_io_clients_0_grant_bits_manager_xact_id ),
       .io_clients_0_grant_bits_is_builtin_type( l1tol2net_io_clients_0_grant_bits_is_builtin_type ),
       .io_clients_0_grant_bits_g_type( l1tol2net_io_clients_0_grant_bits_g_type ),
       .io_clients_0_grant_bits_data( l1tol2net_io_clients_0_grant_bits_data ),
       .io_clients_0_probe_ready( io_tiles_cached_0_probe_ready ),
       .io_clients_0_probe_valid( l1tol2net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_addr_block( l1tol2net_io_clients_0_probe_bits_addr_block ),
       .io_clients_0_probe_bits_p_type( l1tol2net_io_clients_0_probe_bits_p_type ),
       .io_clients_0_release_ready( l1tol2net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_cached_0_release_valid ),
       .io_clients_0_release_bits_addr_beat( io_tiles_cached_0_release_bits_addr_beat ),
       .io_clients_0_release_bits_addr_block( io_tiles_cached_0_release_bits_addr_block ),
       .io_clients_0_release_bits_client_xact_id( io_tiles_cached_0_release_bits_client_xact_id ),
       .io_clients_0_release_bits_r_type( io_tiles_cached_0_release_bits_r_type ),
       .io_clients_0_release_bits_voluntary( io_tiles_cached_0_release_bits_voluntary ),
       .io_clients_0_release_bits_data( io_tiles_cached_0_release_bits_data ),
       .io_managers_0_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_managers_0_acquire_valid( l1tol2net_io_managers_0_acquire_valid ),
       .io_managers_0_acquire_bits_addr_block( l1tol2net_io_managers_0_acquire_bits_addr_block ),
       .io_managers_0_acquire_bits_client_xact_id( l1tol2net_io_managers_0_acquire_bits_client_xact_id ),
       .io_managers_0_acquire_bits_addr_beat( l1tol2net_io_managers_0_acquire_bits_addr_beat ),
       .io_managers_0_acquire_bits_is_builtin_type( l1tol2net_io_managers_0_acquire_bits_is_builtin_type ),
       .io_managers_0_acquire_bits_a_type( l1tol2net_io_managers_0_acquire_bits_a_type ),
       .io_managers_0_acquire_bits_union( l1tol2net_io_managers_0_acquire_bits_union ),
       .io_managers_0_acquire_bits_data( l1tol2net_io_managers_0_acquire_bits_data ),
       .io_managers_0_acquire_bits_client_id( l1tol2net_io_managers_0_acquire_bits_client_id ),
       .io_managers_0_grant_ready( l1tol2net_io_managers_0_grant_ready ),
       .io_managers_0_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_managers_0_grant_bits_addr_beat( L2BroadcastHub_io_inner_grant_bits_addr_beat ),
       .io_managers_0_grant_bits_client_xact_id( L2BroadcastHub_io_inner_grant_bits_client_xact_id ),
       .io_managers_0_grant_bits_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_manager_xact_id ),
       .io_managers_0_grant_bits_is_builtin_type( L2BroadcastHub_io_inner_grant_bits_is_builtin_type ),
       .io_managers_0_grant_bits_g_type( L2BroadcastHub_io_inner_grant_bits_g_type ),
       .io_managers_0_grant_bits_data( L2BroadcastHub_io_inner_grant_bits_data ),
       .io_managers_0_grant_bits_client_id( L2BroadcastHub_io_inner_grant_bits_client_id ),
       .io_managers_0_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_managers_0_finish_valid( l1tol2net_io_managers_0_finish_valid ),
       .io_managers_0_finish_bits_manager_xact_id( l1tol2net_io_managers_0_finish_bits_manager_xact_id ),
       .io_managers_0_probe_ready( l1tol2net_io_managers_0_probe_ready ),
       .io_managers_0_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_managers_0_probe_bits_addr_block( L2BroadcastHub_io_inner_probe_bits_addr_block ),
       .io_managers_0_probe_bits_p_type( L2BroadcastHub_io_inner_probe_bits_p_type ),
       .io_managers_0_probe_bits_client_id( L2BroadcastHub_io_inner_probe_bits_client_id ),
       .io_managers_0_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_managers_0_release_valid( l1tol2net_io_managers_0_release_valid ),
       .io_managers_0_release_bits_addr_beat( l1tol2net_io_managers_0_release_bits_addr_beat ),
       .io_managers_0_release_bits_addr_block( l1tol2net_io_managers_0_release_bits_addr_block ),
       .io_managers_0_release_bits_client_xact_id( l1tol2net_io_managers_0_release_bits_client_xact_id ),
       .io_managers_0_release_bits_r_type( l1tol2net_io_managers_0_release_bits_r_type ),
       .io_managers_0_release_bits_voluntary( l1tol2net_io_managers_0_release_bits_voluntary ),
       .io_managers_0_release_bits_data( l1tol2net_io_managers_0_release_bits_data ),
       .io_managers_0_release_bits_client_id( l1tol2net_io_managers_0_release_bits_client_id )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign l1tol2net.io_clients_2_release_bits_addr_beat = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_addr_block = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_client_xact_id = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_r_type = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_voluntary = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_data = {4{$random}};
    assign l1tol2net.io_clients_1_release_bits_addr_beat = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_addr_block = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_client_xact_id = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_r_type = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_voluntary = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_data = {4{$random}};
// synthesis translate_on
`endif
  L2BroadcastHub L2BroadcastHub(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_inner_acquire_valid( l1tol2net_io_managers_0_acquire_valid ),
       .io_inner_acquire_bits_addr_block( l1tol2net_io_managers_0_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( l1tol2net_io_managers_0_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( l1tol2net_io_managers_0_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( l1tol2net_io_managers_0_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( l1tol2net_io_managers_0_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( l1tol2net_io_managers_0_acquire_bits_union ),
       .io_inner_acquire_bits_data( l1tol2net_io_managers_0_acquire_bits_data ),
       .io_inner_acquire_bits_client_id( l1tol2net_io_managers_0_acquire_bits_client_id ),
       .io_inner_grant_ready( l1tol2net_io_managers_0_grant_ready ),
       .io_inner_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( L2BroadcastHub_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( L2BroadcastHub_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( L2BroadcastHub_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( L2BroadcastHub_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( L2BroadcastHub_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( L2BroadcastHub_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_inner_finish_valid( l1tol2net_io_managers_0_finish_valid ),
       .io_inner_finish_bits_manager_xact_id( l1tol2net_io_managers_0_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( l1tol2net_io_managers_0_probe_ready ),
       .io_inner_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( L2BroadcastHub_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( L2BroadcastHub_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( L2BroadcastHub_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_inner_release_valid( l1tol2net_io_managers_0_release_valid ),
       .io_inner_release_bits_addr_beat( l1tol2net_io_managers_0_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( l1tol2net_io_managers_0_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( l1tol2net_io_managers_0_release_bits_client_xact_id ),
       .io_inner_release_bits_r_type( l1tol2net_io_managers_0_release_bits_r_type ),
       .io_inner_release_bits_voluntary( l1tol2net_io_managers_0_release_bits_voluntary ),
       .io_inner_release_bits_data( l1tol2net_io_managers_0_release_bits_data ),
       .io_inner_release_bits_client_id( l1tol2net_io_managers_0_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( ClientTileLinkIOWrapper_2_io_in_acquire_ready ),
       .io_outer_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( L2BroadcastHub_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( L2BroadcastHub_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( L2BroadcastHub_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( L2BroadcastHub_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( L2BroadcastHub_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( L2BroadcastHub_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_outer_grant_valid( ClientTileLinkIOWrapper_2_io_in_grant_valid ),
       .io_outer_grant_bits_addr_beat( ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type ),
       .io_outer_grant_bits_data( ClientTileLinkIOWrapper_2_io_in_grant_bits_data )
  );
  NastiRecursiveInterconnect_1 interconnect(.clk(clk), .reset(reset),
       .io_masters_1_aw_ready( interconnect_io_masters_1_aw_ready ),
       .io_masters_1_aw_valid( rtc_io_aw_valid ),
       .io_masters_1_aw_bits_addr( rtc_io_aw_bits_addr ),
       .io_masters_1_aw_bits_len( rtc_io_aw_bits_len ),
       .io_masters_1_aw_bits_size( rtc_io_aw_bits_size ),
       .io_masters_1_aw_bits_burst( rtc_io_aw_bits_burst ),
       .io_masters_1_aw_bits_lock( rtc_io_aw_bits_lock ),
       .io_masters_1_aw_bits_cache( rtc_io_aw_bits_cache ),
       .io_masters_1_aw_bits_prot( rtc_io_aw_bits_prot ),
       .io_masters_1_aw_bits_qos( rtc_io_aw_bits_qos ),
       .io_masters_1_aw_bits_region( rtc_io_aw_bits_region ),
       .io_masters_1_aw_bits_id( rtc_io_aw_bits_id ),
       .io_masters_1_aw_bits_user( rtc_io_aw_bits_user ),
       .io_masters_1_w_ready( interconnect_io_masters_1_w_ready ),
       .io_masters_1_w_valid( rtc_io_w_valid ),
       .io_masters_1_w_bits_data( rtc_io_w_bits_data ),
       .io_masters_1_w_bits_last( rtc_io_w_bits_last ),
       .io_masters_1_w_bits_strb( rtc_io_w_bits_strb ),
       .io_masters_1_w_bits_user( rtc_io_w_bits_user ),
       .io_masters_1_b_ready( rtc_io_b_ready ),
       .io_masters_1_b_valid( interconnect_io_masters_1_b_valid ),
       .io_masters_1_b_bits_resp( interconnect_io_masters_1_b_bits_resp ),
       .io_masters_1_b_bits_id( interconnect_io_masters_1_b_bits_id ),
       .io_masters_1_b_bits_user( interconnect_io_masters_1_b_bits_user ),
       .io_masters_1_ar_ready( interconnect_io_masters_1_ar_ready ),
       .io_masters_1_ar_valid( rtc_io_ar_valid ),
       //.io_masters_1_ar_bits_addr(  )
       //.io_masters_1_ar_bits_len(  )
       //.io_masters_1_ar_bits_size(  )
       //.io_masters_1_ar_bits_burst(  )
       //.io_masters_1_ar_bits_lock(  )
       //.io_masters_1_ar_bits_cache(  )
       //.io_masters_1_ar_bits_prot(  )
       //.io_masters_1_ar_bits_qos(  )
       //.io_masters_1_ar_bits_region(  )
       //.io_masters_1_ar_bits_id(  )
       //.io_masters_1_ar_bits_user(  )
       .io_masters_1_r_ready( rtc_io_r_ready ),
       .io_masters_1_r_valid( interconnect_io_masters_1_r_valid ),
       .io_masters_1_r_bits_resp( interconnect_io_masters_1_r_bits_resp ),
       .io_masters_1_r_bits_data( interconnect_io_masters_1_r_bits_data ),
       .io_masters_1_r_bits_last( interconnect_io_masters_1_r_bits_last ),
       .io_masters_1_r_bits_id( interconnect_io_masters_1_r_bits_id ),
       .io_masters_1_r_bits_user( interconnect_io_masters_1_r_bits_user ),
       .io_masters_0_aw_ready( interconnect_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( Queue_1_io_deq_valid ),
       .io_masters_0_aw_bits_addr( Queue_1_io_deq_bits_addr ),
       .io_masters_0_aw_bits_len( Queue_1_io_deq_bits_len ),
       .io_masters_0_aw_bits_size( Queue_1_io_deq_bits_size ),
       .io_masters_0_aw_bits_burst( Queue_1_io_deq_bits_burst ),
       .io_masters_0_aw_bits_lock( Queue_1_io_deq_bits_lock ),
       .io_masters_0_aw_bits_cache( Queue_1_io_deq_bits_cache ),
       .io_masters_0_aw_bits_prot( Queue_1_io_deq_bits_prot ),
       .io_masters_0_aw_bits_qos( Queue_1_io_deq_bits_qos ),
       .io_masters_0_aw_bits_region( Queue_1_io_deq_bits_region ),
       .io_masters_0_aw_bits_id( Queue_1_io_deq_bits_id ),
       .io_masters_0_aw_bits_user( Queue_1_io_deq_bits_user ),
       .io_masters_0_w_ready( interconnect_io_masters_0_w_ready ),
       .io_masters_0_w_valid( Queue_2_io_deq_valid ),
       .io_masters_0_w_bits_data( Queue_2_io_deq_bits_data ),
       .io_masters_0_w_bits_last( Queue_2_io_deq_bits_last ),
       .io_masters_0_w_bits_strb( Queue_2_io_deq_bits_strb ),
       .io_masters_0_w_bits_user( Queue_2_io_deq_bits_user ),
       .io_masters_0_b_ready( Queue_4_io_enq_ready ),
       .io_masters_0_b_valid( interconnect_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( interconnect_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( interconnect_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( interconnect_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( interconnect_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( Queue_io_deq_valid ),
       .io_masters_0_ar_bits_addr( Queue_io_deq_bits_addr ),
       .io_masters_0_ar_bits_len( Queue_io_deq_bits_len ),
       .io_masters_0_ar_bits_size( Queue_io_deq_bits_size ),
       .io_masters_0_ar_bits_burst( Queue_io_deq_bits_burst ),
       .io_masters_0_ar_bits_lock( Queue_io_deq_bits_lock ),
       .io_masters_0_ar_bits_cache( Queue_io_deq_bits_cache ),
       .io_masters_0_ar_bits_prot( Queue_io_deq_bits_prot ),
       .io_masters_0_ar_bits_qos( Queue_io_deq_bits_qos ),
       .io_masters_0_ar_bits_region( Queue_io_deq_bits_region ),
       .io_masters_0_ar_bits_id( Queue_io_deq_bits_id ),
       .io_masters_0_ar_bits_user( Queue_io_deq_bits_user ),
       .io_masters_0_r_ready( Queue_3_io_enq_ready ),
       .io_masters_0_r_valid( interconnect_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( interconnect_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( interconnect_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( interconnect_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( interconnect_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( interconnect_io_masters_0_r_bits_user ),
       .io_slaves_3_aw_ready( io_mmio_aw_ready ),
       .io_slaves_3_aw_valid( interconnect_io_slaves_3_aw_valid ),
       .io_slaves_3_aw_bits_addr( interconnect_io_slaves_3_aw_bits_addr ),
       .io_slaves_3_aw_bits_len( interconnect_io_slaves_3_aw_bits_len ),
       .io_slaves_3_aw_bits_size( interconnect_io_slaves_3_aw_bits_size ),
       .io_slaves_3_aw_bits_burst( interconnect_io_slaves_3_aw_bits_burst ),
       .io_slaves_3_aw_bits_lock( interconnect_io_slaves_3_aw_bits_lock ),
       .io_slaves_3_aw_bits_cache( interconnect_io_slaves_3_aw_bits_cache ),
       .io_slaves_3_aw_bits_prot( interconnect_io_slaves_3_aw_bits_prot ),
       .io_slaves_3_aw_bits_qos( interconnect_io_slaves_3_aw_bits_qos ),
       .io_slaves_3_aw_bits_region( interconnect_io_slaves_3_aw_bits_region ),
       .io_slaves_3_aw_bits_id( interconnect_io_slaves_3_aw_bits_id ),
       .io_slaves_3_aw_bits_user( interconnect_io_slaves_3_aw_bits_user ),
       .io_slaves_3_w_ready( io_mmio_w_ready ),
       .io_slaves_3_w_valid( interconnect_io_slaves_3_w_valid ),
       .io_slaves_3_w_bits_data( interconnect_io_slaves_3_w_bits_data ),
       .io_slaves_3_w_bits_last( interconnect_io_slaves_3_w_bits_last ),
       .io_slaves_3_w_bits_strb( interconnect_io_slaves_3_w_bits_strb ),
       .io_slaves_3_w_bits_user( interconnect_io_slaves_3_w_bits_user ),
       .io_slaves_3_b_ready( interconnect_io_slaves_3_b_ready ),
       .io_slaves_3_b_valid( io_mmio_b_valid ),
       .io_slaves_3_b_bits_resp( io_mmio_b_bits_resp ),
       .io_slaves_3_b_bits_id( io_mmio_b_bits_id ),
       .io_slaves_3_b_bits_user( io_mmio_b_bits_user ),
       .io_slaves_3_ar_ready( io_mmio_ar_ready ),
       .io_slaves_3_ar_valid( interconnect_io_slaves_3_ar_valid ),
       .io_slaves_3_ar_bits_addr( interconnect_io_slaves_3_ar_bits_addr ),
       .io_slaves_3_ar_bits_len( interconnect_io_slaves_3_ar_bits_len ),
       .io_slaves_3_ar_bits_size( interconnect_io_slaves_3_ar_bits_size ),
       .io_slaves_3_ar_bits_burst( interconnect_io_slaves_3_ar_bits_burst ),
       .io_slaves_3_ar_bits_lock( interconnect_io_slaves_3_ar_bits_lock ),
       .io_slaves_3_ar_bits_cache( interconnect_io_slaves_3_ar_bits_cache ),
       .io_slaves_3_ar_bits_prot( interconnect_io_slaves_3_ar_bits_prot ),
       .io_slaves_3_ar_bits_qos( interconnect_io_slaves_3_ar_bits_qos ),
       .io_slaves_3_ar_bits_region( interconnect_io_slaves_3_ar_bits_region ),
       .io_slaves_3_ar_bits_id( interconnect_io_slaves_3_ar_bits_id ),
       .io_slaves_3_ar_bits_user( interconnect_io_slaves_3_ar_bits_user ),
       .io_slaves_3_r_ready( interconnect_io_slaves_3_r_ready ),
       .io_slaves_3_r_valid( io_mmio_r_valid ),
       .io_slaves_3_r_bits_resp( io_mmio_r_bits_resp ),
       .io_slaves_3_r_bits_data( io_mmio_r_bits_data ),
       .io_slaves_3_r_bits_last( io_mmio_r_bits_last ),
       .io_slaves_3_r_bits_id( io_mmio_r_bits_id ),
       .io_slaves_3_r_bits_user( io_mmio_r_bits_user ),
       .io_slaves_2_aw_ready( conv_io_nasti_aw_ready ),
       .io_slaves_2_aw_valid( interconnect_io_slaves_2_aw_valid ),
       .io_slaves_2_aw_bits_addr( interconnect_io_slaves_2_aw_bits_addr ),
       .io_slaves_2_aw_bits_len( interconnect_io_slaves_2_aw_bits_len ),
       .io_slaves_2_aw_bits_size( interconnect_io_slaves_2_aw_bits_size ),
       .io_slaves_2_aw_bits_burst( interconnect_io_slaves_2_aw_bits_burst ),
       .io_slaves_2_aw_bits_lock( interconnect_io_slaves_2_aw_bits_lock ),
       .io_slaves_2_aw_bits_cache( interconnect_io_slaves_2_aw_bits_cache ),
       .io_slaves_2_aw_bits_prot( interconnect_io_slaves_2_aw_bits_prot ),
       .io_slaves_2_aw_bits_qos( interconnect_io_slaves_2_aw_bits_qos ),
       .io_slaves_2_aw_bits_region( interconnect_io_slaves_2_aw_bits_region ),
       .io_slaves_2_aw_bits_id( interconnect_io_slaves_2_aw_bits_id ),
       .io_slaves_2_aw_bits_user( interconnect_io_slaves_2_aw_bits_user ),
       .io_slaves_2_w_ready( conv_io_nasti_w_ready ),
       .io_slaves_2_w_valid( interconnect_io_slaves_2_w_valid ),
       .io_slaves_2_w_bits_data( interconnect_io_slaves_2_w_bits_data ),
       .io_slaves_2_w_bits_last( interconnect_io_slaves_2_w_bits_last ),
       .io_slaves_2_w_bits_strb( interconnect_io_slaves_2_w_bits_strb ),
       .io_slaves_2_w_bits_user( interconnect_io_slaves_2_w_bits_user ),
       .io_slaves_2_b_ready( interconnect_io_slaves_2_b_ready ),
       .io_slaves_2_b_valid( conv_io_nasti_b_valid ),
       .io_slaves_2_b_bits_resp( conv_io_nasti_b_bits_resp ),
       .io_slaves_2_b_bits_id( conv_io_nasti_b_bits_id ),
       .io_slaves_2_b_bits_user( conv_io_nasti_b_bits_user ),
       .io_slaves_2_ar_ready( conv_io_nasti_ar_ready ),
       .io_slaves_2_ar_valid( interconnect_io_slaves_2_ar_valid ),
       .io_slaves_2_ar_bits_addr( interconnect_io_slaves_2_ar_bits_addr ),
       .io_slaves_2_ar_bits_len( interconnect_io_slaves_2_ar_bits_len ),
       .io_slaves_2_ar_bits_size( interconnect_io_slaves_2_ar_bits_size ),
       .io_slaves_2_ar_bits_burst( interconnect_io_slaves_2_ar_bits_burst ),
       .io_slaves_2_ar_bits_lock( interconnect_io_slaves_2_ar_bits_lock ),
       .io_slaves_2_ar_bits_cache( interconnect_io_slaves_2_ar_bits_cache ),
       .io_slaves_2_ar_bits_prot( interconnect_io_slaves_2_ar_bits_prot ),
       .io_slaves_2_ar_bits_qos( interconnect_io_slaves_2_ar_bits_qos ),
       .io_slaves_2_ar_bits_region( interconnect_io_slaves_2_ar_bits_region ),
       .io_slaves_2_ar_bits_id( interconnect_io_slaves_2_ar_bits_id ),
       .io_slaves_2_ar_bits_user( interconnect_io_slaves_2_ar_bits_user ),
       .io_slaves_2_r_ready( interconnect_io_slaves_2_r_ready ),
       .io_slaves_2_r_valid( conv_io_nasti_r_valid ),
       .io_slaves_2_r_bits_resp( conv_io_nasti_r_bits_resp ),
       .io_slaves_2_r_bits_data( conv_io_nasti_r_bits_data ),
       .io_slaves_2_r_bits_last( conv_io_nasti_r_bits_last ),
       .io_slaves_2_r_bits_id( conv_io_nasti_r_bits_id ),
       .io_slaves_2_r_bits_user( conv_io_nasti_r_bits_user ),
       .io_slaves_1_aw_ready( SMIIONastiIOConverter_io_nasti_aw_ready ),
       .io_slaves_1_aw_valid( interconnect_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( interconnect_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( interconnect_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( interconnect_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( interconnect_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( interconnect_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( interconnect_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( interconnect_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( interconnect_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( interconnect_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( interconnect_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( interconnect_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( SMIIONastiIOConverter_io_nasti_w_ready ),
       .io_slaves_1_w_valid( interconnect_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( interconnect_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( interconnect_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( interconnect_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( interconnect_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( interconnect_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( SMIIONastiIOConverter_io_nasti_b_valid ),
       .io_slaves_1_b_bits_resp( SMIIONastiIOConverter_io_nasti_b_bits_resp ),
       .io_slaves_1_b_bits_id( SMIIONastiIOConverter_io_nasti_b_bits_id ),
       .io_slaves_1_b_bits_user( SMIIONastiIOConverter_io_nasti_b_bits_user ),
       .io_slaves_1_ar_ready( SMIIONastiIOConverter_io_nasti_ar_ready ),
       .io_slaves_1_ar_valid( interconnect_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( interconnect_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( interconnect_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( interconnect_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( interconnect_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( interconnect_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( interconnect_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( interconnect_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( interconnect_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( interconnect_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( interconnect_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( interconnect_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( interconnect_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( SMIIONastiIOConverter_io_nasti_r_valid ),
       .io_slaves_1_r_bits_resp( SMIIONastiIOConverter_io_nasti_r_bits_resp ),
       .io_slaves_1_r_bits_data( SMIIONastiIOConverter_io_nasti_r_bits_data ),
       .io_slaves_1_r_bits_last( SMIIONastiIOConverter_io_nasti_r_bits_last ),
       .io_slaves_1_r_bits_id( SMIIONastiIOConverter_io_nasti_r_bits_id ),
       .io_slaves_1_r_bits_user( SMIIONastiIOConverter_io_nasti_r_bits_user ),
       .io_slaves_0_aw_ready( io_mem_0_aw_ready ),
       .io_slaves_0_aw_valid( interconnect_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( interconnect_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( interconnect_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( interconnect_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( interconnect_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( interconnect_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( interconnect_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( interconnect_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( interconnect_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( interconnect_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( interconnect_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( interconnect_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_mem_0_w_ready ),
       .io_slaves_0_w_valid( interconnect_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( interconnect_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( interconnect_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( interconnect_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( interconnect_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( interconnect_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_mem_0_b_valid ),
       .io_slaves_0_b_bits_resp( io_mem_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_mem_0_b_bits_id ),
       .io_slaves_0_b_bits_user( io_mem_0_b_bits_user ),
       .io_slaves_0_ar_ready( io_mem_0_ar_ready ),
       .io_slaves_0_ar_valid( interconnect_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( interconnect_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( interconnect_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( interconnect_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( interconnect_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( interconnect_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( interconnect_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( interconnect_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( interconnect_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( interconnect_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( interconnect_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( interconnect_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( interconnect_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_mem_0_r_valid ),
       .io_slaves_0_r_bits_resp( io_mem_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_mem_0_r_bits_data ),
       .io_slaves_0_r_bits_last( io_mem_0_r_bits_last ),
       .io_slaves_0_r_bits_id( io_mem_0_r_bits_id ),
       .io_slaves_0_r_bits_user( io_mem_0_r_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign interconnect.io_masters_1_ar_bits_addr = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_len = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_size = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_burst = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_lock = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_cache = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_prot = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_qos = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_region = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_id = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_user = {1{$random}};
// synthesis translate_on
`endif
  ClientTileLinkIOUnwrapper ClientTileLinkIOUnwrapper(.clk(clk), .reset(reset),
       .io_in_acquire_ready( ClientTileLinkIOUnwrapper_io_in_acquire_ready ),
       .io_in_acquire_valid( ClientTileLinkIOWrapper_2_io_out_acquire_valid ),
       .io_in_acquire_bits_addr_block( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type ),
       .io_in_acquire_bits_union( ClientTileLinkIOWrapper_2_io_out_acquire_bits_union ),
       .io_in_acquire_bits_data( ClientTileLinkIOWrapper_2_io_out_acquire_bits_data ),
       .io_in_grant_ready( ClientTileLinkIOWrapper_2_io_out_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOUnwrapper_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOUnwrapper_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOUnwrapper_io_in_grant_bits_data ),
       .io_in_probe_ready( ClientTileLinkIOWrapper_2_io_out_probe_ready ),
       .io_in_probe_valid( ClientTileLinkIOUnwrapper_io_in_probe_valid ),
       //.io_in_probe_bits_addr_block(  )
       //.io_in_probe_bits_p_type(  )
       .io_in_release_ready( ClientTileLinkIOUnwrapper_io_in_release_ready ),
       .io_in_release_valid( ClientTileLinkIOWrapper_2_io_out_release_valid ),
       //.io_in_release_bits_addr_beat(  )
       //.io_in_release_bits_addr_block(  )
       //.io_in_release_bits_client_xact_id(  )
       //.io_in_release_bits_r_type(  )
       //.io_in_release_bits_voluntary(  )
       //.io_in_release_bits_data(  )
       .io_out_acquire_ready( TileLinkIONarrower_io_in_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOUnwrapper_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOUnwrapper_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOUnwrapper_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOUnwrapper_io_out_grant_ready ),
       .io_out_grant_valid( TileLinkIONarrower_io_in_grant_valid ),
       .io_out_grant_bits_addr_beat( TileLinkIONarrower_io_in_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( TileLinkIONarrower_io_in_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( TileLinkIONarrower_io_in_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( TileLinkIONarrower_io_in_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( TileLinkIONarrower_io_in_grant_bits_g_type ),
       .io_out_grant_bits_data( TileLinkIONarrower_io_in_grant_bits_data )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ClientTileLinkIOUnwrapper.io_in_release_bits_addr_beat = {1{$random}};
    assign ClientTileLinkIOUnwrapper.io_in_release_bits_addr_block = {1{$random}};
    assign ClientTileLinkIOUnwrapper.io_in_release_bits_client_xact_id = {1{$random}};
    assign ClientTileLinkIOUnwrapper.io_in_release_bits_r_type = {1{$random}};
    assign ClientTileLinkIOUnwrapper.io_in_release_bits_voluntary = {1{$random}};
    assign ClientTileLinkIOUnwrapper.io_in_release_bits_data = {4{$random}};
// synthesis translate_on
`endif
  TileLinkIONarrower TileLinkIONarrower(.clk(clk), .reset(reset),
       .io_in_acquire_ready( TileLinkIONarrower_io_in_acquire_ready ),
       .io_in_acquire_valid( ClientTileLinkIOUnwrapper_io_out_acquire_valid ),
       .io_in_acquire_bits_addr_block( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_out_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_a_type ),
       .io_in_acquire_bits_union( ClientTileLinkIOUnwrapper_io_out_acquire_bits_union ),
       .io_in_acquire_bits_data( ClientTileLinkIOUnwrapper_io_out_acquire_bits_data ),
       .io_in_grant_ready( ClientTileLinkIOUnwrapper_io_out_grant_ready ),
       .io_in_grant_valid( TileLinkIONarrower_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( TileLinkIONarrower_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( TileLinkIONarrower_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( TileLinkIONarrower_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( TileLinkIONarrower_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( TileLinkIONarrower_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( TileLinkIONarrower_io_in_grant_bits_data ),
       .io_out_acquire_ready( NastiIOTileLinkIOConverter_io_tl_acquire_ready ),
       .io_out_acquire_valid( TileLinkIONarrower_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( TileLinkIONarrower_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( TileLinkIONarrower_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( TileLinkIONarrower_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( TileLinkIONarrower_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( TileLinkIONarrower_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( TileLinkIONarrower_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( TileLinkIONarrower_io_out_acquire_bits_data ),
       .io_out_grant_ready( TileLinkIONarrower_io_out_grant_ready ),
       .io_out_grant_valid( NastiIOTileLinkIOConverter_io_tl_grant_valid ),
       .io_out_grant_bits_addr_beat( NastiIOTileLinkIOConverter_io_tl_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_g_type ),
       .io_out_grant_bits_data( NastiIOTileLinkIOConverter_io_tl_grant_bits_data )
  );
  NastiIOTileLinkIOConverter NastiIOTileLinkIOConverter(.clk(clk), .reset(reset),
       .io_tl_acquire_ready( NastiIOTileLinkIOConverter_io_tl_acquire_ready ),
       .io_tl_acquire_valid( TileLinkIONarrower_io_out_acquire_valid ),
       .io_tl_acquire_bits_addr_block( TileLinkIONarrower_io_out_acquire_bits_addr_block ),
       .io_tl_acquire_bits_client_xact_id( TileLinkIONarrower_io_out_acquire_bits_client_xact_id ),
       .io_tl_acquire_bits_addr_beat( TileLinkIONarrower_io_out_acquire_bits_addr_beat ),
       .io_tl_acquire_bits_is_builtin_type( TileLinkIONarrower_io_out_acquire_bits_is_builtin_type ),
       .io_tl_acquire_bits_a_type( TileLinkIONarrower_io_out_acquire_bits_a_type ),
       .io_tl_acquire_bits_union( TileLinkIONarrower_io_out_acquire_bits_union ),
       .io_tl_acquire_bits_data( TileLinkIONarrower_io_out_acquire_bits_data ),
       .io_tl_grant_ready( TileLinkIONarrower_io_out_grant_ready ),
       .io_tl_grant_valid( NastiIOTileLinkIOConverter_io_tl_grant_valid ),
       .io_tl_grant_bits_addr_beat( NastiIOTileLinkIOConverter_io_tl_grant_bits_addr_beat ),
       .io_tl_grant_bits_client_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id ),
       .io_tl_grant_bits_manager_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id ),
       .io_tl_grant_bits_is_builtin_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type ),
       .io_tl_grant_bits_g_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_g_type ),
       .io_tl_grant_bits_data( NastiIOTileLinkIOConverter_io_tl_grant_bits_data ),
       .io_nasti_aw_ready( Queue_1_io_enq_ready ),
       .io_nasti_aw_valid( NastiIOTileLinkIOConverter_io_nasti_aw_valid ),
       .io_nasti_aw_bits_addr( NastiIOTileLinkIOConverter_io_nasti_aw_bits_addr ),
       .io_nasti_aw_bits_len( NastiIOTileLinkIOConverter_io_nasti_aw_bits_len ),
       .io_nasti_aw_bits_size( NastiIOTileLinkIOConverter_io_nasti_aw_bits_size ),
       .io_nasti_aw_bits_burst( NastiIOTileLinkIOConverter_io_nasti_aw_bits_burst ),
       .io_nasti_aw_bits_lock( NastiIOTileLinkIOConverter_io_nasti_aw_bits_lock ),
       .io_nasti_aw_bits_cache( NastiIOTileLinkIOConverter_io_nasti_aw_bits_cache ),
       .io_nasti_aw_bits_prot( NastiIOTileLinkIOConverter_io_nasti_aw_bits_prot ),
       .io_nasti_aw_bits_qos( NastiIOTileLinkIOConverter_io_nasti_aw_bits_qos ),
       .io_nasti_aw_bits_region( NastiIOTileLinkIOConverter_io_nasti_aw_bits_region ),
       .io_nasti_aw_bits_id( NastiIOTileLinkIOConverter_io_nasti_aw_bits_id ),
       .io_nasti_aw_bits_user( NastiIOTileLinkIOConverter_io_nasti_aw_bits_user ),
       .io_nasti_w_ready( Queue_2_io_enq_ready ),
       .io_nasti_w_valid( NastiIOTileLinkIOConverter_io_nasti_w_valid ),
       .io_nasti_w_bits_data( NastiIOTileLinkIOConverter_io_nasti_w_bits_data ),
       .io_nasti_w_bits_last( NastiIOTileLinkIOConverter_io_nasti_w_bits_last ),
       .io_nasti_w_bits_strb( NastiIOTileLinkIOConverter_io_nasti_w_bits_strb ),
       .io_nasti_w_bits_user( NastiIOTileLinkIOConverter_io_nasti_w_bits_user ),
       .io_nasti_b_ready( NastiIOTileLinkIOConverter_io_nasti_b_ready ),
       .io_nasti_b_valid( Queue_4_io_deq_valid ),
       .io_nasti_b_bits_resp( Queue_4_io_deq_bits_resp ),
       .io_nasti_b_bits_id( Queue_4_io_deq_bits_id ),
       .io_nasti_b_bits_user( Queue_4_io_deq_bits_user ),
       .io_nasti_ar_ready( Queue_io_enq_ready ),
       .io_nasti_ar_valid( NastiIOTileLinkIOConverter_io_nasti_ar_valid ),
       .io_nasti_ar_bits_addr( NastiIOTileLinkIOConverter_io_nasti_ar_bits_addr ),
       .io_nasti_ar_bits_len( NastiIOTileLinkIOConverter_io_nasti_ar_bits_len ),
       .io_nasti_ar_bits_size( NastiIOTileLinkIOConverter_io_nasti_ar_bits_size ),
       .io_nasti_ar_bits_burst( NastiIOTileLinkIOConverter_io_nasti_ar_bits_burst ),
       .io_nasti_ar_bits_lock( NastiIOTileLinkIOConverter_io_nasti_ar_bits_lock ),
       .io_nasti_ar_bits_cache( NastiIOTileLinkIOConverter_io_nasti_ar_bits_cache ),
       .io_nasti_ar_bits_prot( NastiIOTileLinkIOConverter_io_nasti_ar_bits_prot ),
       .io_nasti_ar_bits_qos( NastiIOTileLinkIOConverter_io_nasti_ar_bits_qos ),
       .io_nasti_ar_bits_region( NastiIOTileLinkIOConverter_io_nasti_ar_bits_region ),
       .io_nasti_ar_bits_id( NastiIOTileLinkIOConverter_io_nasti_ar_bits_id ),
       .io_nasti_ar_bits_user( NastiIOTileLinkIOConverter_io_nasti_ar_bits_user ),
       .io_nasti_r_ready( NastiIOTileLinkIOConverter_io_nasti_r_ready ),
       .io_nasti_r_valid( Queue_3_io_deq_valid ),
       .io_nasti_r_bits_resp( Queue_3_io_deq_bits_resp ),
       .io_nasti_r_bits_data( Queue_3_io_deq_bits_data ),
       .io_nasti_r_bits_last( Queue_3_io_deq_bits_last ),
       .io_nasti_r_bits_id( Queue_3_io_deq_bits_id ),
       .io_nasti_r_bits_user( Queue_3_io_deq_bits_user )
  );
  ClientTileLinkIOWrapper_1 ClientTileLinkIOWrapper_2(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_2_io_in_acquire_ready ),
       .io_in_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_in_acquire_bits_addr_block( L2BroadcastHub_io_outer_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( L2BroadcastHub_io_outer_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( L2BroadcastHub_io_outer_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( L2BroadcastHub_io_outer_acquire_bits_a_type ),
       .io_in_acquire_bits_union( L2BroadcastHub_io_outer_acquire_bits_union ),
       .io_in_acquire_bits_data( L2BroadcastHub_io_outer_acquire_bits_data ),
       .io_in_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_2_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_2_io_in_grant_bits_data ),
       .io_out_acquire_ready( ClientTileLinkIOUnwrapper_io_in_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_2_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_2_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_2_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_2_io_out_grant_ready ),
       .io_out_grant_valid( ClientTileLinkIOUnwrapper_io_in_grant_valid ),
       .io_out_grant_bits_addr_beat( ClientTileLinkIOUnwrapper_io_in_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_g_type ),
       .io_out_grant_bits_data( ClientTileLinkIOUnwrapper_io_in_grant_bits_data ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_2_io_out_probe_ready ),
       .io_out_probe_valid( ClientTileLinkIOUnwrapper_io_in_probe_valid ),
       //.io_out_probe_bits_addr_block(  )
       //.io_out_probe_bits_p_type(  )
       .io_out_release_ready( ClientTileLinkIOUnwrapper_io_in_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_2_io_out_release_valid )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_data(  )
  );
  Queue_3 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( NastiIOTileLinkIOConverter_io_nasti_ar_valid ),
       .io_enq_bits_addr( NastiIOTileLinkIOConverter_io_nasti_ar_bits_addr ),
       .io_enq_bits_len( NastiIOTileLinkIOConverter_io_nasti_ar_bits_len ),
       .io_enq_bits_size( NastiIOTileLinkIOConverter_io_nasti_ar_bits_size ),
       .io_enq_bits_burst( NastiIOTileLinkIOConverter_io_nasti_ar_bits_burst ),
       .io_enq_bits_lock( NastiIOTileLinkIOConverter_io_nasti_ar_bits_lock ),
       .io_enq_bits_cache( NastiIOTileLinkIOConverter_io_nasti_ar_bits_cache ),
       .io_enq_bits_prot( NastiIOTileLinkIOConverter_io_nasti_ar_bits_prot ),
       .io_enq_bits_qos( NastiIOTileLinkIOConverter_io_nasti_ar_bits_qos ),
       .io_enq_bits_region( NastiIOTileLinkIOConverter_io_nasti_ar_bits_region ),
       .io_enq_bits_id( NastiIOTileLinkIOConverter_io_nasti_ar_bits_id ),
       .io_enq_bits_user( NastiIOTileLinkIOConverter_io_nasti_ar_bits_user ),
       .io_deq_ready( interconnect_io_masters_0_ar_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_io_deq_bits_len ),
       .io_deq_bits_size( Queue_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_io_deq_bits_lock ),
       .io_deq_bits_cache( Queue_io_deq_bits_cache ),
       .io_deq_bits_prot( Queue_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_io_deq_bits_region ),
       .io_deq_bits_id( Queue_io_deq_bits_id ),
       .io_deq_bits_user( Queue_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_3 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( NastiIOTileLinkIOConverter_io_nasti_aw_valid ),
       .io_enq_bits_addr( NastiIOTileLinkIOConverter_io_nasti_aw_bits_addr ),
       .io_enq_bits_len( NastiIOTileLinkIOConverter_io_nasti_aw_bits_len ),
       .io_enq_bits_size( NastiIOTileLinkIOConverter_io_nasti_aw_bits_size ),
       .io_enq_bits_burst( NastiIOTileLinkIOConverter_io_nasti_aw_bits_burst ),
       .io_enq_bits_lock( NastiIOTileLinkIOConverter_io_nasti_aw_bits_lock ),
       .io_enq_bits_cache( NastiIOTileLinkIOConverter_io_nasti_aw_bits_cache ),
       .io_enq_bits_prot( NastiIOTileLinkIOConverter_io_nasti_aw_bits_prot ),
       .io_enq_bits_qos( NastiIOTileLinkIOConverter_io_nasti_aw_bits_qos ),
       .io_enq_bits_region( NastiIOTileLinkIOConverter_io_nasti_aw_bits_region ),
       .io_enq_bits_id( NastiIOTileLinkIOConverter_io_nasti_aw_bits_id ),
       .io_enq_bits_user( NastiIOTileLinkIOConverter_io_nasti_aw_bits_user ),
       .io_deq_ready( interconnect_io_masters_0_aw_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_addr( Queue_1_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_1_io_deq_bits_len ),
       .io_deq_bits_size( Queue_1_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_1_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_1_io_deq_bits_lock ),
       .io_deq_bits_cache( Queue_1_io_deq_bits_cache ),
       .io_deq_bits_prot( Queue_1_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_1_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_1_io_deq_bits_region ),
       .io_deq_bits_id( Queue_1_io_deq_bits_id ),
       .io_deq_bits_user( Queue_1_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_4 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( NastiIOTileLinkIOConverter_io_nasti_w_valid ),
       .io_enq_bits_data( NastiIOTileLinkIOConverter_io_nasti_w_bits_data ),
       .io_enq_bits_last( NastiIOTileLinkIOConverter_io_nasti_w_bits_last ),
       .io_enq_bits_strb( NastiIOTileLinkIOConverter_io_nasti_w_bits_strb ),
       .io_enq_bits_user( NastiIOTileLinkIOConverter_io_nasti_w_bits_user ),
       .io_deq_ready( interconnect_io_masters_0_w_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_data( Queue_2_io_deq_bits_data ),
       .io_deq_bits_last( Queue_2_io_deq_bits_last ),
       .io_deq_bits_strb( Queue_2_io_deq_bits_strb ),
       .io_deq_bits_user( Queue_2_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_5 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( interconnect_io_masters_0_r_valid ),
       .io_enq_bits_resp( interconnect_io_masters_0_r_bits_resp ),
       .io_enq_bits_data( interconnect_io_masters_0_r_bits_data ),
       .io_enq_bits_last( interconnect_io_masters_0_r_bits_last ),
       .io_enq_bits_id( interconnect_io_masters_0_r_bits_id ),
       .io_enq_bits_user( interconnect_io_masters_0_r_bits_user ),
       .io_deq_ready( NastiIOTileLinkIOConverter_io_nasti_r_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_resp( Queue_3_io_deq_bits_resp ),
       .io_deq_bits_data( Queue_3_io_deq_bits_data ),
       .io_deq_bits_last( Queue_3_io_deq_bits_last ),
       .io_deq_bits_id( Queue_3_io_deq_bits_id ),
       .io_deq_bits_user( Queue_3_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_6 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( interconnect_io_masters_0_b_valid ),
       .io_enq_bits_resp( interconnect_io_masters_0_b_bits_resp ),
       .io_enq_bits_id( interconnect_io_masters_0_b_bits_id ),
       .io_enq_bits_user( interconnect_io_masters_0_b_bits_user ),
       .io_deq_ready( NastiIOTileLinkIOConverter_io_nasti_b_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_resp( Queue_4_io_deq_bits_resp ),
       .io_deq_bits_id( Queue_4_io_deq_bits_id ),
       .io_deq_bits_user( Queue_4_io_deq_bits_user )
       //.io_count(  )
  );
  RTC rtc(.clk(clk), .reset(reset),
       .io_aw_ready( interconnect_io_masters_1_aw_ready ),
       .io_aw_valid( rtc_io_aw_valid ),
       .io_aw_bits_addr( rtc_io_aw_bits_addr ),
       .io_aw_bits_len( rtc_io_aw_bits_len ),
       .io_aw_bits_size( rtc_io_aw_bits_size ),
       .io_aw_bits_burst( rtc_io_aw_bits_burst ),
       .io_aw_bits_lock( rtc_io_aw_bits_lock ),
       .io_aw_bits_cache( rtc_io_aw_bits_cache ),
       .io_aw_bits_prot( rtc_io_aw_bits_prot ),
       .io_aw_bits_qos( rtc_io_aw_bits_qos ),
       .io_aw_bits_region( rtc_io_aw_bits_region ),
       .io_aw_bits_id( rtc_io_aw_bits_id ),
       .io_aw_bits_user( rtc_io_aw_bits_user ),
       .io_w_ready( interconnect_io_masters_1_w_ready ),
       .io_w_valid( rtc_io_w_valid ),
       .io_w_bits_data( rtc_io_w_bits_data ),
       .io_w_bits_last( rtc_io_w_bits_last ),
       .io_w_bits_strb( rtc_io_w_bits_strb ),
       .io_w_bits_user( rtc_io_w_bits_user ),
       .io_b_ready( rtc_io_b_ready ),
       .io_b_valid( interconnect_io_masters_1_b_valid ),
       .io_b_bits_resp( interconnect_io_masters_1_b_bits_resp ),
       .io_b_bits_id( interconnect_io_masters_1_b_bits_id ),
       .io_b_bits_user( interconnect_io_masters_1_b_bits_user ),
       .io_ar_ready( interconnect_io_masters_1_ar_ready ),
       .io_ar_valid( rtc_io_ar_valid ),
       //.io_ar_bits_addr(  )
       //.io_ar_bits_len(  )
       //.io_ar_bits_size(  )
       //.io_ar_bits_burst(  )
       //.io_ar_bits_lock(  )
       //.io_ar_bits_cache(  )
       //.io_ar_bits_prot(  )
       //.io_ar_bits_qos(  )
       //.io_ar_bits_region(  )
       //.io_ar_bits_id(  )
       //.io_ar_bits_user(  )
       .io_r_ready( rtc_io_r_ready ),
       .io_r_valid( interconnect_io_masters_1_r_valid ),
       .io_r_bits_resp( interconnect_io_masters_1_r_bits_resp ),
       .io_r_bits_data( interconnect_io_masters_1_r_bits_data ),
       .io_r_bits_last( interconnect_io_masters_1_r_bits_last ),
       .io_r_bits_id( interconnect_io_masters_1_r_bits_id ),
       .io_r_bits_user( interconnect_io_masters_1_r_bits_user )
  );
  SMIIONastiIOConverter_0 SMIIONastiIOConverter(.clk(clk), .reset(reset),
       .io_nasti_aw_ready( SMIIONastiIOConverter_io_nasti_aw_ready ),
       .io_nasti_aw_valid( interconnect_io_slaves_1_aw_valid ),
       .io_nasti_aw_bits_addr( interconnect_io_slaves_1_aw_bits_addr ),
       .io_nasti_aw_bits_len( interconnect_io_slaves_1_aw_bits_len ),
       .io_nasti_aw_bits_size( interconnect_io_slaves_1_aw_bits_size ),
       .io_nasti_aw_bits_burst( interconnect_io_slaves_1_aw_bits_burst ),
       .io_nasti_aw_bits_lock( interconnect_io_slaves_1_aw_bits_lock ),
       .io_nasti_aw_bits_cache( interconnect_io_slaves_1_aw_bits_cache ),
       .io_nasti_aw_bits_prot( interconnect_io_slaves_1_aw_bits_prot ),
       .io_nasti_aw_bits_qos( interconnect_io_slaves_1_aw_bits_qos ),
       .io_nasti_aw_bits_region( interconnect_io_slaves_1_aw_bits_region ),
       .io_nasti_aw_bits_id( interconnect_io_slaves_1_aw_bits_id ),
       .io_nasti_aw_bits_user( interconnect_io_slaves_1_aw_bits_user ),
       .io_nasti_w_ready( SMIIONastiIOConverter_io_nasti_w_ready ),
       .io_nasti_w_valid( interconnect_io_slaves_1_w_valid ),
       .io_nasti_w_bits_data( interconnect_io_slaves_1_w_bits_data ),
       .io_nasti_w_bits_last( interconnect_io_slaves_1_w_bits_last ),
       .io_nasti_w_bits_strb( interconnect_io_slaves_1_w_bits_strb ),
       .io_nasti_w_bits_user( interconnect_io_slaves_1_w_bits_user ),
       .io_nasti_b_ready( interconnect_io_slaves_1_b_ready ),
       .io_nasti_b_valid( SMIIONastiIOConverter_io_nasti_b_valid ),
       .io_nasti_b_bits_resp( SMIIONastiIOConverter_io_nasti_b_bits_resp ),
       .io_nasti_b_bits_id( SMIIONastiIOConverter_io_nasti_b_bits_id ),
       .io_nasti_b_bits_user( SMIIONastiIOConverter_io_nasti_b_bits_user ),
       .io_nasti_ar_ready( SMIIONastiIOConverter_io_nasti_ar_ready ),
       .io_nasti_ar_valid( interconnect_io_slaves_1_ar_valid ),
       .io_nasti_ar_bits_addr( interconnect_io_slaves_1_ar_bits_addr ),
       .io_nasti_ar_bits_len( interconnect_io_slaves_1_ar_bits_len ),
       .io_nasti_ar_bits_size( interconnect_io_slaves_1_ar_bits_size ),
       .io_nasti_ar_bits_burst( interconnect_io_slaves_1_ar_bits_burst ),
       .io_nasti_ar_bits_lock( interconnect_io_slaves_1_ar_bits_lock ),
       .io_nasti_ar_bits_cache( interconnect_io_slaves_1_ar_bits_cache ),
       .io_nasti_ar_bits_prot( interconnect_io_slaves_1_ar_bits_prot ),
       .io_nasti_ar_bits_qos( interconnect_io_slaves_1_ar_bits_qos ),
       .io_nasti_ar_bits_region( interconnect_io_slaves_1_ar_bits_region ),
       .io_nasti_ar_bits_id( interconnect_io_slaves_1_ar_bits_id ),
       .io_nasti_ar_bits_user( interconnect_io_slaves_1_ar_bits_user ),
       .io_nasti_r_ready( interconnect_io_slaves_1_r_ready ),
       .io_nasti_r_valid( SMIIONastiIOConverter_io_nasti_r_valid ),
       .io_nasti_r_bits_resp( SMIIONastiIOConverter_io_nasti_r_bits_resp ),
       .io_nasti_r_bits_data( SMIIONastiIOConverter_io_nasti_r_bits_data ),
       .io_nasti_r_bits_last( SMIIONastiIOConverter_io_nasti_r_bits_last ),
       .io_nasti_r_bits_id( SMIIONastiIOConverter_io_nasti_r_bits_id ),
       .io_nasti_r_bits_user( SMIIONastiIOConverter_io_nasti_r_bits_user ),
       .io_smi_req_ready( io_csr_0_req_ready ),
       .io_smi_req_valid( SMIIONastiIOConverter_io_smi_req_valid ),
       .io_smi_req_bits_rw( SMIIONastiIOConverter_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( SMIIONastiIOConverter_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( SMIIONastiIOConverter_io_smi_req_bits_data ),
       .io_smi_resp_ready( SMIIONastiIOConverter_io_smi_resp_ready ),
       .io_smi_resp_valid( io_csr_0_resp_valid ),
       .io_smi_resp_bits( io_csr_0_resp_bits )
  );
  SMIIONastiIOConverter_1 conv(.clk(clk), .reset(reset),
       .io_nasti_aw_ready( conv_io_nasti_aw_ready ),
       .io_nasti_aw_valid( interconnect_io_slaves_2_aw_valid ),
       .io_nasti_aw_bits_addr( interconnect_io_slaves_2_aw_bits_addr ),
       .io_nasti_aw_bits_len( interconnect_io_slaves_2_aw_bits_len ),
       .io_nasti_aw_bits_size( interconnect_io_slaves_2_aw_bits_size ),
       .io_nasti_aw_bits_burst( interconnect_io_slaves_2_aw_bits_burst ),
       .io_nasti_aw_bits_lock( interconnect_io_slaves_2_aw_bits_lock ),
       .io_nasti_aw_bits_cache( interconnect_io_slaves_2_aw_bits_cache ),
       .io_nasti_aw_bits_prot( interconnect_io_slaves_2_aw_bits_prot ),
       .io_nasti_aw_bits_qos( interconnect_io_slaves_2_aw_bits_qos ),
       .io_nasti_aw_bits_region( interconnect_io_slaves_2_aw_bits_region ),
       .io_nasti_aw_bits_id( interconnect_io_slaves_2_aw_bits_id ),
       .io_nasti_aw_bits_user( interconnect_io_slaves_2_aw_bits_user ),
       .io_nasti_w_ready( conv_io_nasti_w_ready ),
       .io_nasti_w_valid( interconnect_io_slaves_2_w_valid ),
       .io_nasti_w_bits_data( interconnect_io_slaves_2_w_bits_data ),
       .io_nasti_w_bits_last( interconnect_io_slaves_2_w_bits_last ),
       .io_nasti_w_bits_strb( interconnect_io_slaves_2_w_bits_strb ),
       .io_nasti_w_bits_user( interconnect_io_slaves_2_w_bits_user ),
       .io_nasti_b_ready( interconnect_io_slaves_2_b_ready ),
       .io_nasti_b_valid( conv_io_nasti_b_valid ),
       .io_nasti_b_bits_resp( conv_io_nasti_b_bits_resp ),
       .io_nasti_b_bits_id( conv_io_nasti_b_bits_id ),
       .io_nasti_b_bits_user( conv_io_nasti_b_bits_user ),
       .io_nasti_ar_ready( conv_io_nasti_ar_ready ),
       .io_nasti_ar_valid( interconnect_io_slaves_2_ar_valid ),
       .io_nasti_ar_bits_addr( interconnect_io_slaves_2_ar_bits_addr ),
       .io_nasti_ar_bits_len( interconnect_io_slaves_2_ar_bits_len ),
       .io_nasti_ar_bits_size( interconnect_io_slaves_2_ar_bits_size ),
       .io_nasti_ar_bits_burst( interconnect_io_slaves_2_ar_bits_burst ),
       .io_nasti_ar_bits_lock( interconnect_io_slaves_2_ar_bits_lock ),
       .io_nasti_ar_bits_cache( interconnect_io_slaves_2_ar_bits_cache ),
       .io_nasti_ar_bits_prot( interconnect_io_slaves_2_ar_bits_prot ),
       .io_nasti_ar_bits_qos( interconnect_io_slaves_2_ar_bits_qos ),
       .io_nasti_ar_bits_region( interconnect_io_slaves_2_ar_bits_region ),
       .io_nasti_ar_bits_id( interconnect_io_slaves_2_ar_bits_id ),
       .io_nasti_ar_bits_user( interconnect_io_slaves_2_ar_bits_user ),
       .io_nasti_r_ready( interconnect_io_slaves_2_r_ready ),
       .io_nasti_r_valid( conv_io_nasti_r_valid ),
       .io_nasti_r_bits_resp( conv_io_nasti_r_bits_resp ),
       .io_nasti_r_bits_data( conv_io_nasti_r_bits_data ),
       .io_nasti_r_bits_last( conv_io_nasti_r_bits_last ),
       .io_nasti_r_bits_id( conv_io_nasti_r_bits_id ),
       .io_nasti_r_bits_user( conv_io_nasti_r_bits_user ),
       .io_smi_req_ready( io_scr_req_ready ),
       .io_smi_req_valid( conv_io_smi_req_valid ),
       .io_smi_req_bits_rw( conv_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( conv_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( conv_io_smi_req_bits_data ),
       .io_smi_resp_ready( conv_io_smi_resp_ready ),
       .io_smi_resp_valid( io_scr_resp_valid ),
       .io_smi_resp_bits( io_scr_resp_bits )
  );
endmodule

module SCRFile(input clk, input reset,
    output io_smi_req_ready,
    input  io_smi_req_valid,
    input  io_smi_req_bits_rw,
    input [5:0] io_smi_req_bits_addr,
    input [63:0] io_smi_req_bits_data,
    input  io_smi_resp_ready,
    output io_smi_resp_valid,
    output[63:0] io_smi_resp_bits,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    //input [63:0] io_scr_rdata_1
    //input [63:0] io_scr_rdata_0
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[63:0] T5;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T8;
  wire[5:0] T9;
  reg [5:0] read_addr;
  wire[5:0] T135;
  wire[5:0] T10;
  wire T11;
  wire[63:0] T12;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T13;
  wire T14;
  wire[63:0] T15;
  wire[63:0] T16;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T17;
  wire[63:0] T18;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T19;
  wire T20;
  wire T21;
  wire[63:0] T22;
  wire[63:0] T23;
  wire[63:0] T24;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T25;
  wire[63:0] T26;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T27;
  wire T28;
  wire[63:0] T29;
  wire[63:0] T30;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T31;
  wire[63:0] T32;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[63:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T41;
  wire[63:0] T42;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T43;
  wire T44;
  wire[63:0] T45;
  wire[63:0] T46;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T47;
  wire[63:0] T48;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T49;
  wire T50;
  wire T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire[63:0] T54;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T55;
  wire[63:0] T56;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T57;
  wire T58;
  wire[63:0] T59;
  wire[63:0] T60;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T61;
  wire[63:0] T62;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[63:0] T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[63:0] T71;
  wire[63:0] T72;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T73;
  wire[63:0] T74;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T75;
  wire T76;
  wire[63:0] T77;
  wire[63:0] T78;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T79;
  wire[63:0] T80;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T81;
  wire T82;
  wire T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T87;
  wire[63:0] T88;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T89;
  wire T90;
  wire[63:0] T91;
  wire[63:0] T92;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T93;
  wire[63:0] T94;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[63:0] T99;
  wire[63:0] T100;
  wire[63:0] T101;
  wire[63:0] T102;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T103;
  wire[63:0] T104;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T105;
  wire T106;
  wire[63:0] T107;
  wire[63:0] T108;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T109;
  wire[63:0] T110;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T111;
  wire T112;
  wire T113;
  wire[63:0] T114;
  wire[63:0] T115;
  wire[63:0] T116;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T117;
  wire[63:0] T118;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T119;
  wire T120;
  wire[63:0] T121;
  wire[63:0] T122;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T123;
  wire[63:0] T124;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  reg  resp_valid;
  wire T136;
  wire T131;
  wire T132;
  wire T133;
  wire T134;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    read_addr = {1{$random}};
    resp_valid = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_scr_wdata = io_smi_req_bits_data;
  assign io_scr_waddr = io_smi_req_bits_addr;
  assign io_scr_wen = T0;
  assign T0 = T1 & io_smi_req_bits_rw;
  assign T1 = io_smi_req_ready & io_smi_req_valid;
  assign io_smi_resp_bits = T2;
  assign T2 = T130 ? T68 : T3;
  assign T3 = T67 ? T37 : T4;
  assign T4 = T36 ? T22 : T5;
  assign T5 = T21 ? T15 : T6;
  assign T6 = T14 ? T12 : T7;
  assign T7 = T8 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = 64'h1;
  assign scr_rdata_1 = 64'h400;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = read_addr;
  assign T135 = reset ? 6'h0 : T10;
  assign T10 = T11 ? io_smi_req_bits_addr : read_addr;
  assign T11 = io_smi_req_ready & io_smi_req_valid;
  assign T12 = T13 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T13 = T9[1'h0:1'h0];
  assign T14 = T9[1'h1:1'h1];
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign T22 = T35 ? T29 : T23;
  assign T23 = T28 ? T26 : T24;
  assign T24 = T25 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T25 = T9[1'h0:1'h0];
  assign T26 = T27 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T27 = T9[1'h0:1'h0];
  assign T28 = T9[1'h1:1'h1];
  assign T29 = T34 ? T32 : T30;
  assign T30 = T31 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T31 = T9[1'h0:1'h0];
  assign T32 = T33 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T33 = T9[1'h0:1'h0];
  assign T34 = T9[1'h1:1'h1];
  assign T35 = T9[2'h2:2'h2];
  assign T36 = T9[2'h3:2'h3];
  assign T37 = T66 ? T52 : T38;
  assign T38 = T51 ? T45 : T39;
  assign T39 = T44 ? T42 : T40;
  assign T40 = T41 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T41 = T9[1'h0:1'h0];
  assign T42 = T43 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T43 = T9[1'h0:1'h0];
  assign T44 = T9[1'h1:1'h1];
  assign T45 = T50 ? T48 : T46;
  assign T46 = T47 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T47 = T9[1'h0:1'h0];
  assign T48 = T49 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T49 = T9[1'h0:1'h0];
  assign T50 = T9[1'h1:1'h1];
  assign T51 = T9[2'h2:2'h2];
  assign T52 = T65 ? T59 : T53;
  assign T53 = T58 ? T56 : T54;
  assign T54 = T55 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T55 = T9[1'h0:1'h0];
  assign T56 = T57 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T57 = T9[1'h0:1'h0];
  assign T58 = T9[1'h1:1'h1];
  assign T59 = T64 ? T62 : T60;
  assign T60 = T61 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T61 = T9[1'h0:1'h0];
  assign T62 = T63 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T63 = T9[1'h0:1'h0];
  assign T64 = T9[1'h1:1'h1];
  assign T65 = T9[2'h2:2'h2];
  assign T66 = T9[2'h3:2'h3];
  assign T67 = T9[3'h4:3'h4];
  assign T68 = T129 ? T99 : T69;
  assign T69 = T98 ? T84 : T70;
  assign T70 = T83 ? T77 : T71;
  assign T71 = T76 ? T74 : T72;
  assign T72 = T73 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T73 = T9[1'h0:1'h0];
  assign T74 = T75 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T75 = T9[1'h0:1'h0];
  assign T76 = T9[1'h1:1'h1];
  assign T77 = T82 ? T80 : T78;
  assign T78 = T79 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T79 = T9[1'h0:1'h0];
  assign T80 = T81 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T81 = T9[1'h0:1'h0];
  assign T82 = T9[1'h1:1'h1];
  assign T83 = T9[2'h2:2'h2];
  assign T84 = T97 ? T91 : T85;
  assign T85 = T90 ? T88 : T86;
  assign T86 = T87 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T87 = T9[1'h0:1'h0];
  assign T88 = T89 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T89 = T9[1'h0:1'h0];
  assign T90 = T9[1'h1:1'h1];
  assign T91 = T96 ? T94 : T92;
  assign T92 = T93 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T93 = T9[1'h0:1'h0];
  assign T94 = T95 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T95 = T9[1'h0:1'h0];
  assign T96 = T9[1'h1:1'h1];
  assign T97 = T9[2'h2:2'h2];
  assign T98 = T9[2'h3:2'h3];
  assign T99 = T128 ? T114 : T100;
  assign T100 = T113 ? T107 : T101;
  assign T101 = T106 ? T104 : T102;
  assign T102 = T103 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T103 = T9[1'h0:1'h0];
  assign T104 = T105 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T105 = T9[1'h0:1'h0];
  assign T106 = T9[1'h1:1'h1];
  assign T107 = T112 ? T110 : T108;
  assign T108 = T109 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T109 = T9[1'h0:1'h0];
  assign T110 = T111 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T111 = T9[1'h0:1'h0];
  assign T112 = T9[1'h1:1'h1];
  assign T113 = T9[2'h2:2'h2];
  assign T114 = T127 ? T121 : T115;
  assign T115 = T120 ? T118 : T116;
  assign T116 = T117 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T117 = T9[1'h0:1'h0];
  assign T118 = T119 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T119 = T9[1'h0:1'h0];
  assign T120 = T9[1'h1:1'h1];
  assign T121 = T126 ? T124 : T122;
  assign T122 = T123 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T123 = T9[1'h0:1'h0];
  assign T124 = T125 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T125 = T9[1'h0:1'h0];
  assign T126 = T9[1'h1:1'h1];
  assign T127 = T9[2'h2:2'h2];
  assign T128 = T9[2'h3:2'h3];
  assign T129 = T9[3'h4:3'h4];
  assign T130 = T9[3'h5:3'h5];
  assign io_smi_resp_valid = resp_valid;
  assign T136 = reset ? 1'h0 : T131;
  assign T131 = T133 ? 1'h0 : T132;
  assign T132 = T11 ? 1'h1 : resp_valid;
  assign T133 = io_smi_resp_ready & io_smi_resp_valid;
  assign io_smi_req_ready = T134;
  assign T134 = resp_valid ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      read_addr <= 6'h0;
    end else if(T11) begin
      read_addr <= io_smi_req_bits_addr;
    end
    if(reset) begin
      resp_valid <= 1'h0;
    end else if(T133) begin
      resp_valid <= 1'h0;
    end else if(T11) begin
      resp_valid <= 1'h1;
    end
  end
endmodule

module Uncore(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_csr,
    input  io_mem_0_aw_ready,
    output io_mem_0_aw_valid,
    output[31:0] io_mem_0_aw_bits_addr,
    output[7:0] io_mem_0_aw_bits_len,
    output[2:0] io_mem_0_aw_bits_size,
    output[1:0] io_mem_0_aw_bits_burst,
    output io_mem_0_aw_bits_lock,
    output[3:0] io_mem_0_aw_bits_cache,
    output[2:0] io_mem_0_aw_bits_prot,
    output[3:0] io_mem_0_aw_bits_qos,
    output[3:0] io_mem_0_aw_bits_region,
    output[4:0] io_mem_0_aw_bits_id,
    output io_mem_0_aw_bits_user,
    input  io_mem_0_w_ready,
    output io_mem_0_w_valid,
    output[63:0] io_mem_0_w_bits_data,
    output io_mem_0_w_bits_last,
    output[7:0] io_mem_0_w_bits_strb,
    output io_mem_0_w_bits_user,
    output io_mem_0_b_ready,
    input  io_mem_0_b_valid,
    input [1:0] io_mem_0_b_bits_resp,
    input [4:0] io_mem_0_b_bits_id,
    input  io_mem_0_b_bits_user,
    input  io_mem_0_ar_ready,
    output io_mem_0_ar_valid,
    output[31:0] io_mem_0_ar_bits_addr,
    output[7:0] io_mem_0_ar_bits_len,
    output[2:0] io_mem_0_ar_bits_size,
    output[1:0] io_mem_0_ar_bits_burst,
    output io_mem_0_ar_bits_lock,
    output[3:0] io_mem_0_ar_bits_cache,
    output[2:0] io_mem_0_ar_bits_prot,
    output[3:0] io_mem_0_ar_bits_qos,
    output[3:0] io_mem_0_ar_bits_region,
    output[4:0] io_mem_0_ar_bits_id,
    output io_mem_0_ar_bits_user,
    output io_mem_0_r_ready,
    input  io_mem_0_r_valid,
    input [1:0] io_mem_0_r_bits_resp,
    input [63:0] io_mem_0_r_bits_data,
    input  io_mem_0_r_bits_last,
    input [4:0] io_mem_0_r_bits_id,
    input  io_mem_0_r_bits_user,
    output io_tiles_cached_0_acquire_ready,
    input  io_tiles_cached_0_acquire_valid,
    input [25:0] io_tiles_cached_0_acquire_bits_addr_block,
    input [1:0] io_tiles_cached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_acquire_bits_addr_beat,
    input  io_tiles_cached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_cached_0_acquire_bits_a_type,
    input [16:0] io_tiles_cached_0_acquire_bits_union,
    input [127:0] io_tiles_cached_0_acquire_bits_data,
    input  io_tiles_cached_0_grant_ready,
    output io_tiles_cached_0_grant_valid,
    output[1:0] io_tiles_cached_0_grant_bits_addr_beat,
    output[1:0] io_tiles_cached_0_grant_bits_client_xact_id,
    output[3:0] io_tiles_cached_0_grant_bits_manager_xact_id,
    output io_tiles_cached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_cached_0_grant_bits_g_type,
    output[127:0] io_tiles_cached_0_grant_bits_data,
    input  io_tiles_cached_0_probe_ready,
    output io_tiles_cached_0_probe_valid,
    output[25:0] io_tiles_cached_0_probe_bits_addr_block,
    output[1:0] io_tiles_cached_0_probe_bits_p_type,
    output io_tiles_cached_0_release_ready,
    input  io_tiles_cached_0_release_valid,
    input [1:0] io_tiles_cached_0_release_bits_addr_beat,
    input [25:0] io_tiles_cached_0_release_bits_addr_block,
    input [1:0] io_tiles_cached_0_release_bits_client_xact_id,
    input [2:0] io_tiles_cached_0_release_bits_r_type,
    input  io_tiles_cached_0_release_bits_voluntary,
    input [127:0] io_tiles_cached_0_release_bits_data,
    output io_tiles_uncached_0_acquire_ready,
    input  io_tiles_uncached_0_acquire_valid,
    input [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
    input [1:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_uncached_0_acquire_bits_addr_beat,
    input  io_tiles_uncached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_uncached_0_acquire_bits_a_type,
    input [16:0] io_tiles_uncached_0_acquire_bits_union,
    input [127:0] io_tiles_uncached_0_acquire_bits_data,
    input  io_tiles_uncached_0_grant_ready,
    output io_tiles_uncached_0_grant_valid,
    output[1:0] io_tiles_uncached_0_grant_bits_addr_beat,
    output[1:0] io_tiles_uncached_0_grant_bits_client_xact_id,
    output[3:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
    output io_tiles_uncached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_uncached_0_grant_bits_g_type,
    output[127:0] io_tiles_uncached_0_grant_bits_data,
    output io_htif_0_reset,
    output io_htif_0_id,
    input  io_htif_0_csr_req_ready,
    output io_htif_0_csr_req_valid,
    output io_htif_0_csr_req_bits_rw,
    output[11:0] io_htif_0_csr_req_bits_addr,
    output[63:0] io_htif_0_csr_req_bits_data,
    output io_htif_0_csr_resp_ready,
    input  io_htif_0_csr_resp_valid,
    input [63:0] io_htif_0_csr_resp_bits,
    output io_htif_0_ipi_req_ready,
    input  io_htif_0_ipi_req_valid,
    input  io_htif_0_ipi_req_bits,
    input  io_htif_0_ipi_rep_ready,
    output io_htif_0_ipi_rep_valid,
    output io_htif_0_ipi_rep_bits,
    input  io_htif_0_debug_stats_csr,
    //input  io_mem_backup_ctrl_en
    //input  io_mem_backup_ctrl_in_valid
    //input  io_mem_backup_ctrl_out_ready
    //output io_mem_backup_ctrl_out_valid
    input  io_mmio_aw_ready,
    output io_mmio_aw_valid,
    output[31:0] io_mmio_aw_bits_addr,
    output[7:0] io_mmio_aw_bits_len,
    output[2:0] io_mmio_aw_bits_size,
    output[1:0] io_mmio_aw_bits_burst,
    output io_mmio_aw_bits_lock,
    output[3:0] io_mmio_aw_bits_cache,
    output[2:0] io_mmio_aw_bits_prot,
    output[3:0] io_mmio_aw_bits_qos,
    output[3:0] io_mmio_aw_bits_region,
    output[4:0] io_mmio_aw_bits_id,
    output io_mmio_aw_bits_user,
    input  io_mmio_w_ready,
    output io_mmio_w_valid,
    output[63:0] io_mmio_w_bits_data,
    output io_mmio_w_bits_last,
    output[7:0] io_mmio_w_bits_strb,
    output io_mmio_w_bits_user,
    output io_mmio_b_ready,
    input  io_mmio_b_valid,
    input [1:0] io_mmio_b_bits_resp,
    input [4:0] io_mmio_b_bits_id,
    input  io_mmio_b_bits_user,
    input  io_mmio_ar_ready,
    output io_mmio_ar_valid,
    output[31:0] io_mmio_ar_bits_addr,
    output[7:0] io_mmio_ar_bits_len,
    output[2:0] io_mmio_ar_bits_size,
    output[1:0] io_mmio_ar_bits_burst,
    output io_mmio_ar_bits_lock,
    output[3:0] io_mmio_ar_bits_cache,
    output[2:0] io_mmio_ar_bits_prot,
    output[3:0] io_mmio_ar_bits_qos,
    output[3:0] io_mmio_ar_bits_region,
    output[4:0] io_mmio_ar_bits_id,
    output io_mmio_ar_bits_user,
    output io_mmio_r_ready,
    input  io_mmio_r_valid,
    input [1:0] io_mmio_r_bits_resp,
    input [63:0] io_mmio_r_bits_data,
    input  io_mmio_r_bits_last,
    input [4:0] io_mmio_r_bits_id,
    input  io_mmio_r_bits_user
);

  wire htif_io_host_in_ready;
  wire htif_io_host_out_valid;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_debug_stats_csr;
  wire htif_io_cpu_0_reset;
  wire htif_io_cpu_0_id;
  wire htif_io_cpu_0_csr_req_valid;
  wire htif_io_cpu_0_csr_req_bits_rw;
  wire[11:0] htif_io_cpu_0_csr_req_bits_addr;
  wire[63:0] htif_io_cpu_0_csr_req_bits_data;
  wire htif_io_cpu_0_csr_resp_ready;
  wire htif_io_cpu_0_ipi_req_ready;
  wire htif_io_cpu_0_ipi_rep_valid;
  wire htif_io_mem_acquire_valid;
  wire[25:0] htif_io_mem_acquire_bits_addr_block;
  wire[1:0] htif_io_mem_acquire_bits_client_xact_id;
  wire[1:0] htif_io_mem_acquire_bits_addr_beat;
  wire htif_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] htif_io_mem_acquire_bits_a_type;
  wire[16:0] htif_io_mem_acquire_bits_union;
  wire[127:0] htif_io_mem_acquire_bits_data;
  wire htif_io_mem_grant_ready;
  wire htif_io_scr_req_valid;
  wire htif_io_scr_req_bits_rw;
  wire[5:0] htif_io_scr_req_bits_addr;
  wire[63:0] htif_io_scr_req_bits_data;
  wire htif_io_scr_resp_ready;
  wire scrFile_io_smi_req_ready;
  wire scrFile_io_smi_resp_valid;
  wire[63:0] scrFile_io_smi_resp_bits;
  wire SMIArbiter_io_in_1_req_ready;
  wire SMIArbiter_io_in_1_resp_valid;
  wire[63:0] SMIArbiter_io_in_1_resp_bits;
  wire SMIArbiter_io_in_0_req_ready;
  wire SMIArbiter_io_in_0_resp_valid;
  wire[63:0] SMIArbiter_io_in_0_resp_bits;
  wire SMIArbiter_io_out_req_valid;
  wire SMIArbiter_io_out_req_bits_rw;
  wire[11:0] SMIArbiter_io_out_req_bits_addr;
  wire[63:0] SMIArbiter_io_out_req_bits_data;
  wire SMIArbiter_io_out_resp_ready;
  wire scrArb_io_in_1_req_ready;
  wire scrArb_io_in_1_resp_valid;
  wire[63:0] scrArb_io_in_1_resp_bits;
  wire scrArb_io_in_0_req_ready;
  wire scrArb_io_in_0_resp_valid;
  wire[63:0] scrArb_io_in_0_resp_bits;
  wire scrArb_io_out_req_valid;
  wire scrArb_io_out_req_bits_rw;
  wire[5:0] scrArb_io_out_req_bits_addr;
  wire[63:0] scrArb_io_out_req_bits_data;
  wire scrArb_io_out_resp_ready;
  wire outmemsys_io_tiles_cached_0_acquire_ready;
  wire outmemsys_io_tiles_cached_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  wire[1:0] outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  wire[3:0] outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_tiles_cached_0_grant_bits_g_type;
  wire[127:0] outmemsys_io_tiles_cached_0_grant_bits_data;
  wire outmemsys_io_tiles_cached_0_probe_valid;
  wire[25:0] outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  wire[1:0] outmemsys_io_tiles_cached_0_probe_bits_p_type;
  wire outmemsys_io_tiles_cached_0_release_ready;
  wire outmemsys_io_tiles_uncached_0_acquire_ready;
  wire outmemsys_io_tiles_uncached_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  wire[1:0] outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire[3:0] outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  wire[127:0] outmemsys_io_tiles_uncached_0_grant_bits_data;
  wire outmemsys_io_htif_uncached_acquire_ready;
  wire outmemsys_io_htif_uncached_grant_valid;
  wire[1:0] outmemsys_io_htif_uncached_grant_bits_addr_beat;
  wire[1:0] outmemsys_io_htif_uncached_grant_bits_client_xact_id;
  wire[3:0] outmemsys_io_htif_uncached_grant_bits_manager_xact_id;
  wire outmemsys_io_htif_uncached_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_htif_uncached_grant_bits_g_type;
  wire[127:0] outmemsys_io_htif_uncached_grant_bits_data;
  wire outmemsys_io_mem_0_aw_valid;
  wire[31:0] outmemsys_io_mem_0_aw_bits_addr;
  wire[7:0] outmemsys_io_mem_0_aw_bits_len;
  wire[2:0] outmemsys_io_mem_0_aw_bits_size;
  wire[1:0] outmemsys_io_mem_0_aw_bits_burst;
  wire outmemsys_io_mem_0_aw_bits_lock;
  wire[3:0] outmemsys_io_mem_0_aw_bits_cache;
  wire[2:0] outmemsys_io_mem_0_aw_bits_prot;
  wire[3:0] outmemsys_io_mem_0_aw_bits_qos;
  wire[3:0] outmemsys_io_mem_0_aw_bits_region;
  wire[4:0] outmemsys_io_mem_0_aw_bits_id;
  wire outmemsys_io_mem_0_aw_bits_user;
  wire outmemsys_io_mem_0_w_valid;
  wire[63:0] outmemsys_io_mem_0_w_bits_data;
  wire outmemsys_io_mem_0_w_bits_last;
  wire[7:0] outmemsys_io_mem_0_w_bits_strb;
  wire outmemsys_io_mem_0_w_bits_user;
  wire outmemsys_io_mem_0_b_ready;
  wire outmemsys_io_mem_0_ar_valid;
  wire[31:0] outmemsys_io_mem_0_ar_bits_addr;
  wire[7:0] outmemsys_io_mem_0_ar_bits_len;
  wire[2:0] outmemsys_io_mem_0_ar_bits_size;
  wire[1:0] outmemsys_io_mem_0_ar_bits_burst;
  wire outmemsys_io_mem_0_ar_bits_lock;
  wire[3:0] outmemsys_io_mem_0_ar_bits_cache;
  wire[2:0] outmemsys_io_mem_0_ar_bits_prot;
  wire[3:0] outmemsys_io_mem_0_ar_bits_qos;
  wire[3:0] outmemsys_io_mem_0_ar_bits_region;
  wire[4:0] outmemsys_io_mem_0_ar_bits_id;
  wire outmemsys_io_mem_0_ar_bits_user;
  wire outmemsys_io_mem_0_r_ready;
  wire outmemsys_io_csr_0_req_valid;
  wire outmemsys_io_csr_0_req_bits_rw;
  wire[11:0] outmemsys_io_csr_0_req_bits_addr;
  wire[63:0] outmemsys_io_csr_0_req_bits_data;
  wire outmemsys_io_csr_0_resp_ready;
  wire outmemsys_io_scr_req_valid;
  wire outmemsys_io_scr_req_bits_rw;
  wire[5:0] outmemsys_io_scr_req_bits_addr;
  wire[63:0] outmemsys_io_scr_req_bits_data;
  wire outmemsys_io_scr_resp_ready;
  wire outmemsys_io_mmio_aw_valid;
  wire[31:0] outmemsys_io_mmio_aw_bits_addr;
  wire[7:0] outmemsys_io_mmio_aw_bits_len;
  wire[2:0] outmemsys_io_mmio_aw_bits_size;
  wire[1:0] outmemsys_io_mmio_aw_bits_burst;
  wire outmemsys_io_mmio_aw_bits_lock;
  wire[3:0] outmemsys_io_mmio_aw_bits_cache;
  wire[2:0] outmemsys_io_mmio_aw_bits_prot;
  wire[3:0] outmemsys_io_mmio_aw_bits_qos;
  wire[3:0] outmemsys_io_mmio_aw_bits_region;
  wire[4:0] outmemsys_io_mmio_aw_bits_id;
  wire outmemsys_io_mmio_aw_bits_user;
  wire outmemsys_io_mmio_w_valid;
  wire[63:0] outmemsys_io_mmio_w_bits_data;
  wire outmemsys_io_mmio_w_bits_last;
  wire[7:0] outmemsys_io_mmio_w_bits_strb;
  wire outmemsys_io_mmio_w_bits_user;
  wire outmemsys_io_mmio_b_ready;
  wire outmemsys_io_mmio_ar_valid;
  wire[31:0] outmemsys_io_mmio_ar_bits_addr;
  wire[7:0] outmemsys_io_mmio_ar_bits_len;
  wire[2:0] outmemsys_io_mmio_ar_bits_size;
  wire[1:0] outmemsys_io_mmio_ar_bits_burst;
  wire outmemsys_io_mmio_ar_bits_lock;
  wire[3:0] outmemsys_io_mmio_ar_bits_cache;
  wire[2:0] outmemsys_io_mmio_ar_bits_prot;
  wire[3:0] outmemsys_io_mmio_ar_bits_qos;
  wire[3:0] outmemsys_io_mmio_ar_bits_region;
  wire[4:0] outmemsys_io_mmio_ar_bits_id;
  wire outmemsys_io_mmio_ar_bits_user;
  wire outmemsys_io_mmio_r_ready;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_backup_ctrl_out_valid = {1{$random}};
  assign io_htif_0_ipi_rep_bits = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign io_mmio_r_ready = outmemsys_io_mmio_r_ready;
  assign io_mmio_ar_bits_user = outmemsys_io_mmio_ar_bits_user;
  assign io_mmio_ar_bits_id = outmemsys_io_mmio_ar_bits_id;
  assign io_mmio_ar_bits_region = outmemsys_io_mmio_ar_bits_region;
  assign io_mmio_ar_bits_qos = outmemsys_io_mmio_ar_bits_qos;
  assign io_mmio_ar_bits_prot = outmemsys_io_mmio_ar_bits_prot;
  assign io_mmio_ar_bits_cache = outmemsys_io_mmio_ar_bits_cache;
  assign io_mmio_ar_bits_lock = outmemsys_io_mmio_ar_bits_lock;
  assign io_mmio_ar_bits_burst = outmemsys_io_mmio_ar_bits_burst;
  assign io_mmio_ar_bits_size = outmemsys_io_mmio_ar_bits_size;
  assign io_mmio_ar_bits_len = outmemsys_io_mmio_ar_bits_len;
  assign io_mmio_ar_bits_addr = outmemsys_io_mmio_ar_bits_addr;
  assign io_mmio_ar_valid = outmemsys_io_mmio_ar_valid;
  assign io_mmio_b_ready = outmemsys_io_mmio_b_ready;
  assign io_mmio_w_bits_user = outmemsys_io_mmio_w_bits_user;
  assign io_mmio_w_bits_strb = outmemsys_io_mmio_w_bits_strb;
  assign io_mmio_w_bits_last = outmemsys_io_mmio_w_bits_last;
  assign io_mmio_w_bits_data = outmemsys_io_mmio_w_bits_data;
  assign io_mmio_w_valid = outmemsys_io_mmio_w_valid;
  assign io_mmio_aw_bits_user = outmemsys_io_mmio_aw_bits_user;
  assign io_mmio_aw_bits_id = outmemsys_io_mmio_aw_bits_id;
  assign io_mmio_aw_bits_region = outmemsys_io_mmio_aw_bits_region;
  assign io_mmio_aw_bits_qos = outmemsys_io_mmio_aw_bits_qos;
  assign io_mmio_aw_bits_prot = outmemsys_io_mmio_aw_bits_prot;
  assign io_mmio_aw_bits_cache = outmemsys_io_mmio_aw_bits_cache;
  assign io_mmio_aw_bits_lock = outmemsys_io_mmio_aw_bits_lock;
  assign io_mmio_aw_bits_burst = outmemsys_io_mmio_aw_bits_burst;
  assign io_mmio_aw_bits_size = outmemsys_io_mmio_aw_bits_size;
  assign io_mmio_aw_bits_len = outmemsys_io_mmio_aw_bits_len;
  assign io_mmio_aw_bits_addr = outmemsys_io_mmio_aw_bits_addr;
  assign io_mmio_aw_valid = outmemsys_io_mmio_aw_valid;
  assign io_htif_0_ipi_rep_valid = htif_io_cpu_0_ipi_rep_valid;
  assign io_htif_0_ipi_req_ready = htif_io_cpu_0_ipi_req_ready;
  assign io_htif_0_csr_resp_ready = SMIArbiter_io_out_resp_ready;
  assign io_htif_0_csr_req_bits_data = SMIArbiter_io_out_req_bits_data;
  assign io_htif_0_csr_req_bits_addr = SMIArbiter_io_out_req_bits_addr;
  assign io_htif_0_csr_req_bits_rw = SMIArbiter_io_out_req_bits_rw;
  assign io_htif_0_csr_req_valid = SMIArbiter_io_out_req_valid;
  assign io_htif_0_id = htif_io_cpu_0_id;
  assign io_tiles_uncached_0_grant_bits_data = outmemsys_io_tiles_uncached_0_grant_bits_data;
  assign io_tiles_uncached_0_grant_bits_g_type = outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_addr_beat = outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_valid = outmemsys_io_tiles_uncached_0_grant_valid;
  assign io_tiles_uncached_0_acquire_ready = outmemsys_io_tiles_uncached_0_acquire_ready;
  assign io_tiles_cached_0_release_ready = outmemsys_io_tiles_cached_0_release_ready;
  assign io_tiles_cached_0_probe_bits_p_type = outmemsys_io_tiles_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_probe_bits_addr_block = outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_valid = outmemsys_io_tiles_cached_0_probe_valid;
  assign io_tiles_cached_0_grant_bits_data = outmemsys_io_tiles_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_g_type = outmemsys_io_tiles_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_client_xact_id = outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_addr_beat = outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_valid = outmemsys_io_tiles_cached_0_grant_valid;
  assign io_tiles_cached_0_acquire_ready = outmemsys_io_tiles_cached_0_acquire_ready;
  assign io_mem_0_r_ready = outmemsys_io_mem_0_r_ready;
  assign io_mem_0_ar_bits_user = outmemsys_io_mem_0_ar_bits_user;
  assign io_mem_0_ar_bits_id = outmemsys_io_mem_0_ar_bits_id;
  assign io_mem_0_ar_bits_region = outmemsys_io_mem_0_ar_bits_region;
  assign io_mem_0_ar_bits_qos = outmemsys_io_mem_0_ar_bits_qos;
  assign io_mem_0_ar_bits_prot = outmemsys_io_mem_0_ar_bits_prot;
  assign io_mem_0_ar_bits_cache = outmemsys_io_mem_0_ar_bits_cache;
  assign io_mem_0_ar_bits_lock = outmemsys_io_mem_0_ar_bits_lock;
  assign io_mem_0_ar_bits_burst = outmemsys_io_mem_0_ar_bits_burst;
  assign io_mem_0_ar_bits_size = outmemsys_io_mem_0_ar_bits_size;
  assign io_mem_0_ar_bits_len = outmemsys_io_mem_0_ar_bits_len;
  assign io_mem_0_ar_bits_addr = outmemsys_io_mem_0_ar_bits_addr;
  assign io_mem_0_ar_valid = outmemsys_io_mem_0_ar_valid;
  assign io_mem_0_b_ready = outmemsys_io_mem_0_b_ready;
  assign io_mem_0_w_bits_user = outmemsys_io_mem_0_w_bits_user;
  assign io_mem_0_w_bits_strb = outmemsys_io_mem_0_w_bits_strb;
  assign io_mem_0_w_bits_last = outmemsys_io_mem_0_w_bits_last;
  assign io_mem_0_w_bits_data = outmemsys_io_mem_0_w_bits_data;
  assign io_mem_0_w_valid = outmemsys_io_mem_0_w_valid;
  assign io_mem_0_aw_bits_user = outmemsys_io_mem_0_aw_bits_user;
  assign io_mem_0_aw_bits_id = outmemsys_io_mem_0_aw_bits_id;
  assign io_mem_0_aw_bits_region = outmemsys_io_mem_0_aw_bits_region;
  assign io_mem_0_aw_bits_qos = outmemsys_io_mem_0_aw_bits_qos;
  assign io_mem_0_aw_bits_prot = outmemsys_io_mem_0_aw_bits_prot;
  assign io_mem_0_aw_bits_cache = outmemsys_io_mem_0_aw_bits_cache;
  assign io_mem_0_aw_bits_lock = outmemsys_io_mem_0_aw_bits_lock;
  assign io_mem_0_aw_bits_burst = outmemsys_io_mem_0_aw_bits_burst;
  assign io_mem_0_aw_bits_size = outmemsys_io_mem_0_aw_bits_size;
  assign io_mem_0_aw_bits_len = outmemsys_io_mem_0_aw_bits_len;
  assign io_mem_0_aw_bits_addr = outmemsys_io_mem_0_aw_bits_addr;
  assign io_mem_0_aw_valid = outmemsys_io_mem_0_aw_valid;
  assign io_host_debug_stats_csr = htif_io_host_debug_stats_csr;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_in_ready = htif_io_host_in_ready;
  Htif htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       .io_host_debug_stats_csr( htif_io_host_debug_stats_csr ),
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       .io_cpu_0_id( htif_io_cpu_0_id ),
       .io_cpu_0_csr_req_ready( SMIArbiter_io_in_0_req_ready ),
       .io_cpu_0_csr_req_valid( htif_io_cpu_0_csr_req_valid ),
       .io_cpu_0_csr_req_bits_rw( htif_io_cpu_0_csr_req_bits_rw ),
       .io_cpu_0_csr_req_bits_addr( htif_io_cpu_0_csr_req_bits_addr ),
       .io_cpu_0_csr_req_bits_data( htif_io_cpu_0_csr_req_bits_data ),
       .io_cpu_0_csr_resp_ready( htif_io_cpu_0_csr_resp_ready ),
       .io_cpu_0_csr_resp_valid( SMIArbiter_io_in_0_resp_valid ),
       .io_cpu_0_csr_resp_bits( SMIArbiter_io_in_0_resp_bits ),
       .io_cpu_0_ipi_req_ready( htif_io_cpu_0_ipi_req_ready ),
       .io_cpu_0_ipi_req_valid( io_htif_0_ipi_req_valid ),
       .io_cpu_0_ipi_req_bits( io_htif_0_ipi_req_bits ),
       .io_cpu_0_ipi_rep_ready( io_htif_0_ipi_rep_ready ),
       .io_cpu_0_ipi_rep_valid( htif_io_cpu_0_ipi_rep_valid ),
       //.io_cpu_0_ipi_rep_bits(  )
       .io_cpu_0_debug_stats_csr( io_htif_0_debug_stats_csr ),
       .io_mem_acquire_ready( outmemsys_io_htif_uncached_acquire_ready ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( htif_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( htif_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( htif_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( htif_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( htif_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( htif_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( htif_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( outmemsys_io_htif_uncached_grant_valid ),
       .io_mem_grant_bits_addr_beat( outmemsys_io_htif_uncached_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( outmemsys_io_htif_uncached_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( outmemsys_io_htif_uncached_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( outmemsys_io_htif_uncached_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( outmemsys_io_htif_uncached_grant_bits_g_type ),
       .io_mem_grant_bits_data( outmemsys_io_htif_uncached_grant_bits_data ),
       .io_scr_req_ready( scrArb_io_in_0_req_ready ),
       .io_scr_req_valid( htif_io_scr_req_valid ),
       .io_scr_req_bits_rw( htif_io_scr_req_bits_rw ),
       .io_scr_req_bits_addr( htif_io_scr_req_bits_addr ),
       .io_scr_req_bits_data( htif_io_scr_req_bits_data ),
       .io_scr_resp_ready( htif_io_scr_resp_ready ),
       .io_scr_resp_valid( scrArb_io_in_0_resp_valid ),
       .io_scr_resp_bits( scrArb_io_in_0_resp_bits )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign htif.io_cpu_0_id = {1{$random}};
// synthesis translate_on
`endif
  OuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_cached_0_acquire_ready( outmemsys_io_tiles_cached_0_acquire_ready ),
       .io_tiles_cached_0_acquire_valid( io_tiles_cached_0_acquire_valid ),
       .io_tiles_cached_0_acquire_bits_addr_block( io_tiles_cached_0_acquire_bits_addr_block ),
       .io_tiles_cached_0_acquire_bits_client_xact_id( io_tiles_cached_0_acquire_bits_client_xact_id ),
       .io_tiles_cached_0_acquire_bits_addr_beat( io_tiles_cached_0_acquire_bits_addr_beat ),
       .io_tiles_cached_0_acquire_bits_is_builtin_type( io_tiles_cached_0_acquire_bits_is_builtin_type ),
       .io_tiles_cached_0_acquire_bits_a_type( io_tiles_cached_0_acquire_bits_a_type ),
       .io_tiles_cached_0_acquire_bits_union( io_tiles_cached_0_acquire_bits_union ),
       .io_tiles_cached_0_acquire_bits_data( io_tiles_cached_0_acquire_bits_data ),
       .io_tiles_cached_0_grant_ready( io_tiles_cached_0_grant_ready ),
       .io_tiles_cached_0_grant_valid( outmemsys_io_tiles_cached_0_grant_valid ),
       .io_tiles_cached_0_grant_bits_addr_beat( outmemsys_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_tiles_cached_0_grant_bits_client_xact_id( outmemsys_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_tiles_cached_0_grant_bits_manager_xact_id( outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_tiles_cached_0_grant_bits_is_builtin_type( outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_tiles_cached_0_grant_bits_g_type( outmemsys_io_tiles_cached_0_grant_bits_g_type ),
       .io_tiles_cached_0_grant_bits_data( outmemsys_io_tiles_cached_0_grant_bits_data ),
       .io_tiles_cached_0_probe_ready( io_tiles_cached_0_probe_ready ),
       .io_tiles_cached_0_probe_valid( outmemsys_io_tiles_cached_0_probe_valid ),
       .io_tiles_cached_0_probe_bits_addr_block( outmemsys_io_tiles_cached_0_probe_bits_addr_block ),
       .io_tiles_cached_0_probe_bits_p_type( outmemsys_io_tiles_cached_0_probe_bits_p_type ),
       .io_tiles_cached_0_release_ready( outmemsys_io_tiles_cached_0_release_ready ),
       .io_tiles_cached_0_release_valid( io_tiles_cached_0_release_valid ),
       .io_tiles_cached_0_release_bits_addr_beat( io_tiles_cached_0_release_bits_addr_beat ),
       .io_tiles_cached_0_release_bits_addr_block( io_tiles_cached_0_release_bits_addr_block ),
       .io_tiles_cached_0_release_bits_client_xact_id( io_tiles_cached_0_release_bits_client_xact_id ),
       .io_tiles_cached_0_release_bits_r_type( io_tiles_cached_0_release_bits_r_type ),
       .io_tiles_cached_0_release_bits_voluntary( io_tiles_cached_0_release_bits_voluntary ),
       .io_tiles_cached_0_release_bits_data( io_tiles_cached_0_release_bits_data ),
       .io_tiles_uncached_0_acquire_ready( outmemsys_io_tiles_uncached_0_acquire_ready ),
       .io_tiles_uncached_0_acquire_valid( io_tiles_uncached_0_acquire_valid ),
       .io_tiles_uncached_0_acquire_bits_addr_block( io_tiles_uncached_0_acquire_bits_addr_block ),
       .io_tiles_uncached_0_acquire_bits_client_xact_id( io_tiles_uncached_0_acquire_bits_client_xact_id ),
       .io_tiles_uncached_0_acquire_bits_addr_beat( io_tiles_uncached_0_acquire_bits_addr_beat ),
       .io_tiles_uncached_0_acquire_bits_is_builtin_type( io_tiles_uncached_0_acquire_bits_is_builtin_type ),
       .io_tiles_uncached_0_acquire_bits_a_type( io_tiles_uncached_0_acquire_bits_a_type ),
       .io_tiles_uncached_0_acquire_bits_union( io_tiles_uncached_0_acquire_bits_union ),
       .io_tiles_uncached_0_acquire_bits_data( io_tiles_uncached_0_acquire_bits_data ),
       .io_tiles_uncached_0_grant_ready( io_tiles_uncached_0_grant_ready ),
       .io_tiles_uncached_0_grant_valid( outmemsys_io_tiles_uncached_0_grant_valid ),
       .io_tiles_uncached_0_grant_bits_addr_beat( outmemsys_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_tiles_uncached_0_grant_bits_client_xact_id( outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_tiles_uncached_0_grant_bits_manager_xact_id( outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_tiles_uncached_0_grant_bits_is_builtin_type( outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_tiles_uncached_0_grant_bits_g_type( outmemsys_io_tiles_uncached_0_grant_bits_g_type ),
       .io_tiles_uncached_0_grant_bits_data( outmemsys_io_tiles_uncached_0_grant_bits_data ),
       .io_htif_uncached_acquire_ready( outmemsys_io_htif_uncached_acquire_ready ),
       .io_htif_uncached_acquire_valid( htif_io_mem_acquire_valid ),
       .io_htif_uncached_acquire_bits_addr_block( htif_io_mem_acquire_bits_addr_block ),
       .io_htif_uncached_acquire_bits_client_xact_id( htif_io_mem_acquire_bits_client_xact_id ),
       .io_htif_uncached_acquire_bits_addr_beat( htif_io_mem_acquire_bits_addr_beat ),
       .io_htif_uncached_acquire_bits_is_builtin_type( htif_io_mem_acquire_bits_is_builtin_type ),
       .io_htif_uncached_acquire_bits_a_type( htif_io_mem_acquire_bits_a_type ),
       .io_htif_uncached_acquire_bits_union( htif_io_mem_acquire_bits_union ),
       .io_htif_uncached_acquire_bits_data( htif_io_mem_acquire_bits_data ),
       .io_htif_uncached_grant_ready( htif_io_mem_grant_ready ),
       .io_htif_uncached_grant_valid( outmemsys_io_htif_uncached_grant_valid ),
       .io_htif_uncached_grant_bits_addr_beat( outmemsys_io_htif_uncached_grant_bits_addr_beat ),
       .io_htif_uncached_grant_bits_client_xact_id( outmemsys_io_htif_uncached_grant_bits_client_xact_id ),
       .io_htif_uncached_grant_bits_manager_xact_id( outmemsys_io_htif_uncached_grant_bits_manager_xact_id ),
       .io_htif_uncached_grant_bits_is_builtin_type( outmemsys_io_htif_uncached_grant_bits_is_builtin_type ),
       .io_htif_uncached_grant_bits_g_type( outmemsys_io_htif_uncached_grant_bits_g_type ),
       .io_htif_uncached_grant_bits_data( outmemsys_io_htif_uncached_grant_bits_data ),
       .io_incoherent_0( htif_io_cpu_0_reset ),
       .io_mem_0_aw_ready( io_mem_0_aw_ready ),
       .io_mem_0_aw_valid( outmemsys_io_mem_0_aw_valid ),
       .io_mem_0_aw_bits_addr( outmemsys_io_mem_0_aw_bits_addr ),
       .io_mem_0_aw_bits_len( outmemsys_io_mem_0_aw_bits_len ),
       .io_mem_0_aw_bits_size( outmemsys_io_mem_0_aw_bits_size ),
       .io_mem_0_aw_bits_burst( outmemsys_io_mem_0_aw_bits_burst ),
       .io_mem_0_aw_bits_lock( outmemsys_io_mem_0_aw_bits_lock ),
       .io_mem_0_aw_bits_cache( outmemsys_io_mem_0_aw_bits_cache ),
       .io_mem_0_aw_bits_prot( outmemsys_io_mem_0_aw_bits_prot ),
       .io_mem_0_aw_bits_qos( outmemsys_io_mem_0_aw_bits_qos ),
       .io_mem_0_aw_bits_region( outmemsys_io_mem_0_aw_bits_region ),
       .io_mem_0_aw_bits_id( outmemsys_io_mem_0_aw_bits_id ),
       .io_mem_0_aw_bits_user( outmemsys_io_mem_0_aw_bits_user ),
       .io_mem_0_w_ready( io_mem_0_w_ready ),
       .io_mem_0_w_valid( outmemsys_io_mem_0_w_valid ),
       .io_mem_0_w_bits_data( outmemsys_io_mem_0_w_bits_data ),
       .io_mem_0_w_bits_last( outmemsys_io_mem_0_w_bits_last ),
       .io_mem_0_w_bits_strb( outmemsys_io_mem_0_w_bits_strb ),
       .io_mem_0_w_bits_user( outmemsys_io_mem_0_w_bits_user ),
       .io_mem_0_b_ready( outmemsys_io_mem_0_b_ready ),
       .io_mem_0_b_valid( io_mem_0_b_valid ),
       .io_mem_0_b_bits_resp( io_mem_0_b_bits_resp ),
       .io_mem_0_b_bits_id( io_mem_0_b_bits_id ),
       .io_mem_0_b_bits_user( io_mem_0_b_bits_user ),
       .io_mem_0_ar_ready( io_mem_0_ar_ready ),
       .io_mem_0_ar_valid( outmemsys_io_mem_0_ar_valid ),
       .io_mem_0_ar_bits_addr( outmemsys_io_mem_0_ar_bits_addr ),
       .io_mem_0_ar_bits_len( outmemsys_io_mem_0_ar_bits_len ),
       .io_mem_0_ar_bits_size( outmemsys_io_mem_0_ar_bits_size ),
       .io_mem_0_ar_bits_burst( outmemsys_io_mem_0_ar_bits_burst ),
       .io_mem_0_ar_bits_lock( outmemsys_io_mem_0_ar_bits_lock ),
       .io_mem_0_ar_bits_cache( outmemsys_io_mem_0_ar_bits_cache ),
       .io_mem_0_ar_bits_prot( outmemsys_io_mem_0_ar_bits_prot ),
       .io_mem_0_ar_bits_qos( outmemsys_io_mem_0_ar_bits_qos ),
       .io_mem_0_ar_bits_region( outmemsys_io_mem_0_ar_bits_region ),
       .io_mem_0_ar_bits_id( outmemsys_io_mem_0_ar_bits_id ),
       .io_mem_0_ar_bits_user( outmemsys_io_mem_0_ar_bits_user ),
       .io_mem_0_r_ready( outmemsys_io_mem_0_r_ready ),
       .io_mem_0_r_valid( io_mem_0_r_valid ),
       .io_mem_0_r_bits_resp( io_mem_0_r_bits_resp ),
       .io_mem_0_r_bits_data( io_mem_0_r_bits_data ),
       .io_mem_0_r_bits_last( io_mem_0_r_bits_last ),
       .io_mem_0_r_bits_id( io_mem_0_r_bits_id ),
       .io_mem_0_r_bits_user( io_mem_0_r_bits_user ),
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
       .io_csr_0_req_ready( SMIArbiter_io_in_1_req_ready ),
       .io_csr_0_req_valid( outmemsys_io_csr_0_req_valid ),
       .io_csr_0_req_bits_rw( outmemsys_io_csr_0_req_bits_rw ),
       .io_csr_0_req_bits_addr( outmemsys_io_csr_0_req_bits_addr ),
       .io_csr_0_req_bits_data( outmemsys_io_csr_0_req_bits_data ),
       .io_csr_0_resp_ready( outmemsys_io_csr_0_resp_ready ),
       .io_csr_0_resp_valid( SMIArbiter_io_in_1_resp_valid ),
       .io_csr_0_resp_bits( SMIArbiter_io_in_1_resp_bits ),
       .io_scr_req_ready( scrArb_io_in_1_req_ready ),
       .io_scr_req_valid( outmemsys_io_scr_req_valid ),
       .io_scr_req_bits_rw( outmemsys_io_scr_req_bits_rw ),
       .io_scr_req_bits_addr( outmemsys_io_scr_req_bits_addr ),
       .io_scr_req_bits_data( outmemsys_io_scr_req_bits_data ),
       .io_scr_resp_ready( outmemsys_io_scr_resp_ready ),
       .io_scr_resp_valid( scrArb_io_in_1_resp_valid ),
       .io_scr_resp_bits( scrArb_io_in_1_resp_bits ),
       .io_mmio_aw_ready( io_mmio_aw_ready ),
       .io_mmio_aw_valid( outmemsys_io_mmio_aw_valid ),
       .io_mmio_aw_bits_addr( outmemsys_io_mmio_aw_bits_addr ),
       .io_mmio_aw_bits_len( outmemsys_io_mmio_aw_bits_len ),
       .io_mmio_aw_bits_size( outmemsys_io_mmio_aw_bits_size ),
       .io_mmio_aw_bits_burst( outmemsys_io_mmio_aw_bits_burst ),
       .io_mmio_aw_bits_lock( outmemsys_io_mmio_aw_bits_lock ),
       .io_mmio_aw_bits_cache( outmemsys_io_mmio_aw_bits_cache ),
       .io_mmio_aw_bits_prot( outmemsys_io_mmio_aw_bits_prot ),
       .io_mmio_aw_bits_qos( outmemsys_io_mmio_aw_bits_qos ),
       .io_mmio_aw_bits_region( outmemsys_io_mmio_aw_bits_region ),
       .io_mmio_aw_bits_id( outmemsys_io_mmio_aw_bits_id ),
       .io_mmio_aw_bits_user( outmemsys_io_mmio_aw_bits_user ),
       .io_mmio_w_ready( io_mmio_w_ready ),
       .io_mmio_w_valid( outmemsys_io_mmio_w_valid ),
       .io_mmio_w_bits_data( outmemsys_io_mmio_w_bits_data ),
       .io_mmio_w_bits_last( outmemsys_io_mmio_w_bits_last ),
       .io_mmio_w_bits_strb( outmemsys_io_mmio_w_bits_strb ),
       .io_mmio_w_bits_user( outmemsys_io_mmio_w_bits_user ),
       .io_mmio_b_ready( outmemsys_io_mmio_b_ready ),
       .io_mmio_b_valid( io_mmio_b_valid ),
       .io_mmio_b_bits_resp( io_mmio_b_bits_resp ),
       .io_mmio_b_bits_id( io_mmio_b_bits_id ),
       .io_mmio_b_bits_user( io_mmio_b_bits_user ),
       .io_mmio_ar_ready( io_mmio_ar_ready ),
       .io_mmio_ar_valid( outmemsys_io_mmio_ar_valid ),
       .io_mmio_ar_bits_addr( outmemsys_io_mmio_ar_bits_addr ),
       .io_mmio_ar_bits_len( outmemsys_io_mmio_ar_bits_len ),
       .io_mmio_ar_bits_size( outmemsys_io_mmio_ar_bits_size ),
       .io_mmio_ar_bits_burst( outmemsys_io_mmio_ar_bits_burst ),
       .io_mmio_ar_bits_lock( outmemsys_io_mmio_ar_bits_lock ),
       .io_mmio_ar_bits_cache( outmemsys_io_mmio_ar_bits_cache ),
       .io_mmio_ar_bits_prot( outmemsys_io_mmio_ar_bits_prot ),
       .io_mmio_ar_bits_qos( outmemsys_io_mmio_ar_bits_qos ),
       .io_mmio_ar_bits_region( outmemsys_io_mmio_ar_bits_region ),
       .io_mmio_ar_bits_id( outmemsys_io_mmio_ar_bits_id ),
       .io_mmio_ar_bits_user( outmemsys_io_mmio_ar_bits_user ),
       .io_mmio_r_ready( outmemsys_io_mmio_r_ready ),
       .io_mmio_r_valid( io_mmio_r_valid ),
       .io_mmio_r_bits_resp( io_mmio_r_bits_resp ),
       .io_mmio_r_bits_data( io_mmio_r_bits_data ),
       .io_mmio_r_bits_last( io_mmio_r_bits_last ),
       .io_mmio_r_bits_id( io_mmio_r_bits_id ),
       .io_mmio_r_bits_user( io_mmio_r_bits_user )
  );
  SMIArbiter_0 SMIArbiter(.clk(clk), .reset(reset),
       .io_in_1_req_ready( SMIArbiter_io_in_1_req_ready ),
       .io_in_1_req_valid( outmemsys_io_csr_0_req_valid ),
       .io_in_1_req_bits_rw( outmemsys_io_csr_0_req_bits_rw ),
       .io_in_1_req_bits_addr( outmemsys_io_csr_0_req_bits_addr ),
       .io_in_1_req_bits_data( outmemsys_io_csr_0_req_bits_data ),
       .io_in_1_resp_ready( outmemsys_io_csr_0_resp_ready ),
       .io_in_1_resp_valid( SMIArbiter_io_in_1_resp_valid ),
       .io_in_1_resp_bits( SMIArbiter_io_in_1_resp_bits ),
       .io_in_0_req_ready( SMIArbiter_io_in_0_req_ready ),
       .io_in_0_req_valid( htif_io_cpu_0_csr_req_valid ),
       .io_in_0_req_bits_rw( htif_io_cpu_0_csr_req_bits_rw ),
       .io_in_0_req_bits_addr( htif_io_cpu_0_csr_req_bits_addr ),
       .io_in_0_req_bits_data( htif_io_cpu_0_csr_req_bits_data ),
       .io_in_0_resp_ready( htif_io_cpu_0_csr_resp_ready ),
       .io_in_0_resp_valid( SMIArbiter_io_in_0_resp_valid ),
       .io_in_0_resp_bits( SMIArbiter_io_in_0_resp_bits ),
       .io_out_req_ready( io_htif_0_csr_req_ready ),
       .io_out_req_valid( SMIArbiter_io_out_req_valid ),
       .io_out_req_bits_rw( SMIArbiter_io_out_req_bits_rw ),
       .io_out_req_bits_addr( SMIArbiter_io_out_req_bits_addr ),
       .io_out_req_bits_data( SMIArbiter_io_out_req_bits_data ),
       .io_out_resp_ready( SMIArbiter_io_out_resp_ready ),
       .io_out_resp_valid( io_htif_0_csr_resp_valid ),
       .io_out_resp_bits( io_htif_0_csr_resp_bits )
  );
  SCRFile scrFile(.clk(clk), .reset(reset),
       .io_smi_req_ready( scrFile_io_smi_req_ready ),
       .io_smi_req_valid( scrArb_io_out_req_valid ),
       .io_smi_req_bits_rw( scrArb_io_out_req_bits_rw ),
       .io_smi_req_bits_addr( scrArb_io_out_req_bits_addr ),
       .io_smi_req_bits_data( scrArb_io_out_req_bits_data ),
       .io_smi_resp_ready( scrArb_io_out_resp_ready ),
       .io_smi_resp_valid( scrFile_io_smi_resp_valid ),
       .io_smi_resp_bits( scrFile_io_smi_resp_bits )
       //.io_scr_rdata_63(  )
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       //.io_scr_rdata_2(  )
       //.io_scr_rdata_1(  )
       //.io_scr_rdata_0(  )
       //.io_scr_wen(  )
       //.io_scr_waddr(  )
       //.io_scr_wdata(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign scrFile.io_scr_rdata_63 = {2{$random}};
    assign scrFile.io_scr_rdata_62 = {2{$random}};
    assign scrFile.io_scr_rdata_61 = {2{$random}};
    assign scrFile.io_scr_rdata_60 = {2{$random}};
    assign scrFile.io_scr_rdata_59 = {2{$random}};
    assign scrFile.io_scr_rdata_58 = {2{$random}};
    assign scrFile.io_scr_rdata_57 = {2{$random}};
    assign scrFile.io_scr_rdata_56 = {2{$random}};
    assign scrFile.io_scr_rdata_55 = {2{$random}};
    assign scrFile.io_scr_rdata_54 = {2{$random}};
    assign scrFile.io_scr_rdata_53 = {2{$random}};
    assign scrFile.io_scr_rdata_52 = {2{$random}};
    assign scrFile.io_scr_rdata_51 = {2{$random}};
    assign scrFile.io_scr_rdata_50 = {2{$random}};
    assign scrFile.io_scr_rdata_49 = {2{$random}};
    assign scrFile.io_scr_rdata_48 = {2{$random}};
    assign scrFile.io_scr_rdata_47 = {2{$random}};
    assign scrFile.io_scr_rdata_46 = {2{$random}};
    assign scrFile.io_scr_rdata_45 = {2{$random}};
    assign scrFile.io_scr_rdata_44 = {2{$random}};
    assign scrFile.io_scr_rdata_43 = {2{$random}};
    assign scrFile.io_scr_rdata_42 = {2{$random}};
    assign scrFile.io_scr_rdata_41 = {2{$random}};
    assign scrFile.io_scr_rdata_40 = {2{$random}};
    assign scrFile.io_scr_rdata_39 = {2{$random}};
    assign scrFile.io_scr_rdata_38 = {2{$random}};
    assign scrFile.io_scr_rdata_37 = {2{$random}};
    assign scrFile.io_scr_rdata_36 = {2{$random}};
    assign scrFile.io_scr_rdata_35 = {2{$random}};
    assign scrFile.io_scr_rdata_34 = {2{$random}};
    assign scrFile.io_scr_rdata_33 = {2{$random}};
    assign scrFile.io_scr_rdata_32 = {2{$random}};
    assign scrFile.io_scr_rdata_31 = {2{$random}};
    assign scrFile.io_scr_rdata_30 = {2{$random}};
    assign scrFile.io_scr_rdata_29 = {2{$random}};
    assign scrFile.io_scr_rdata_28 = {2{$random}};
    assign scrFile.io_scr_rdata_27 = {2{$random}};
    assign scrFile.io_scr_rdata_26 = {2{$random}};
    assign scrFile.io_scr_rdata_25 = {2{$random}};
    assign scrFile.io_scr_rdata_24 = {2{$random}};
    assign scrFile.io_scr_rdata_23 = {2{$random}};
    assign scrFile.io_scr_rdata_22 = {2{$random}};
    assign scrFile.io_scr_rdata_21 = {2{$random}};
    assign scrFile.io_scr_rdata_20 = {2{$random}};
    assign scrFile.io_scr_rdata_19 = {2{$random}};
    assign scrFile.io_scr_rdata_18 = {2{$random}};
    assign scrFile.io_scr_rdata_17 = {2{$random}};
    assign scrFile.io_scr_rdata_16 = {2{$random}};
    assign scrFile.io_scr_rdata_15 = {2{$random}};
    assign scrFile.io_scr_rdata_14 = {2{$random}};
    assign scrFile.io_scr_rdata_13 = {2{$random}};
    assign scrFile.io_scr_rdata_12 = {2{$random}};
    assign scrFile.io_scr_rdata_11 = {2{$random}};
    assign scrFile.io_scr_rdata_10 = {2{$random}};
    assign scrFile.io_scr_rdata_9 = {2{$random}};
    assign scrFile.io_scr_rdata_8 = {2{$random}};
    assign scrFile.io_scr_rdata_7 = {2{$random}};
    assign scrFile.io_scr_rdata_6 = {2{$random}};
    assign scrFile.io_scr_rdata_5 = {2{$random}};
    assign scrFile.io_scr_rdata_4 = {2{$random}};
    assign scrFile.io_scr_rdata_3 = {2{$random}};
    assign scrFile.io_scr_rdata_2 = {2{$random}};
// synthesis translate_on
`endif
  SMIArbiter_1 scrArb(.clk(clk), .reset(reset),
       .io_in_1_req_ready( scrArb_io_in_1_req_ready ),
       .io_in_1_req_valid( outmemsys_io_scr_req_valid ),
       .io_in_1_req_bits_rw( outmemsys_io_scr_req_bits_rw ),
       .io_in_1_req_bits_addr( outmemsys_io_scr_req_bits_addr ),
       .io_in_1_req_bits_data( outmemsys_io_scr_req_bits_data ),
       .io_in_1_resp_ready( outmemsys_io_scr_resp_ready ),
       .io_in_1_resp_valid( scrArb_io_in_1_resp_valid ),
       .io_in_1_resp_bits( scrArb_io_in_1_resp_bits ),
       .io_in_0_req_ready( scrArb_io_in_0_req_ready ),
       .io_in_0_req_valid( htif_io_scr_req_valid ),
       .io_in_0_req_bits_rw( htif_io_scr_req_bits_rw ),
       .io_in_0_req_bits_addr( htif_io_scr_req_bits_addr ),
       .io_in_0_req_bits_data( htif_io_scr_req_bits_data ),
       .io_in_0_resp_ready( htif_io_scr_resp_ready ),
       .io_in_0_resp_valid( scrArb_io_in_0_resp_valid ),
       .io_in_0_resp_bits( scrArb_io_in_0_resp_bits ),
       .io_out_req_ready( scrFile_io_smi_req_ready ),
       .io_out_req_valid( scrArb_io_out_req_valid ),
       .io_out_req_bits_rw( scrArb_io_out_req_bits_rw ),
       .io_out_req_bits_addr( scrArb_io_out_req_bits_addr ),
       .io_out_req_bits_data( scrArb_io_out_req_bits_data ),
       .io_out_resp_ready( scrArb_io_out_resp_ready ),
       .io_out_resp_valid( scrFile_io_smi_resp_valid ),
       .io_out_resp_bits( scrFile_io_smi_resp_bits )
  );
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_csr_req_ready,
    input  io_host_csr_req_valid,
    input  io_host_csr_req_bits_rw,
    input [11:0] io_host_csr_req_bits_addr,
    input [63:0] io_host_csr_req_bits_data,
    input  io_host_csr_resp_ready,
    output io_host_csr_resp_valid,
    output[63:0] io_host_csr_resp_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_csr,
    input [11:0] io_rw_addr,
    input [2:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    output io_csr_replay,
    output io_csr_stall,
    output io_csr_xcpt,
    output io_eret,
    output io_status_sd,
    output[30:0] io_status_zero2,
    output io_status_sd_rv32,
    output[8:0] io_status_zero1,
    output[4:0] io_status_vm,
    output io_status_mprv,
    output[1:0] io_status_xs,
    output[1:0] io_status_fs,
    output[1:0] io_status_prv3,
    output io_status_ie3,
    output[1:0] io_status_prv2,
    output io_status_ie2,
    output[1:0] io_status_prv1,
    output io_status_ie1,
    output[1:0] io_status_prv,
    output io_status_ie,
    output[31:0] io_ptbr,
    output[39:0] io_evec,
    input  io_exception,
    input  io_retire,
    input  io_uarch_counters_15,
    input  io_uarch_counters_14,
    input  io_uarch_counters_13,
    input  io_uarch_counters_12,
    input  io_uarch_counters_11,
    input  io_uarch_counters_10,
    input  io_uarch_counters_9,
    input  io_uarch_counters_8,
    input  io_uarch_counters_7,
    input  io_uarch_counters_6,
    input  io_uarch_counters_5,
    input  io_uarch_counters_4,
    input  io_uarch_counters_3,
    input  io_uarch_counters_2,
    input  io_uarch_counters_1,
    input  io_uarch_counters_0,
    input [63:0] io_cause,
    input [39:0] io_pc,
    output io_fatc,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input [39:0] io_rocc_mem_req_bits_addr,
    input [8:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_kill,
    input  io_rocc_mem_req_bits_phys,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[39:0] io_rocc_mem_resp_bits_addr
    //output[8:0] io_rocc_mem_resp_bits_tag
    //output[4:0] io_rocc_mem_resp_bits_cmd
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_word_bypass
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[8:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_invalidate_lr,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [25:0] io_rocc_imem_acquire_bits_addr_block,
    input [1:0] io_rocc_imem_acquire_bits_client_xact_id,
    input [1:0] io_rocc_imem_acquire_bits_addr_beat,
    input  io_rocc_imem_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_imem_acquire_bits_a_type,
    input [16:0] io_rocc_imem_acquire_bits_union,
    input [127:0] io_rocc_imem_acquire_bits_data,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_addr_beat
    //output[1:0] io_rocc_imem_grant_bits_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_manager_xact_id
    //output io_rocc_imem_grant_bits_is_builtin_type
    //output[3:0] io_rocc_imem_grant_bits_g_type
    //output[127:0] io_rocc_imem_grant_bits_data
    //output io_rocc_dmem_0_acquire_ready
    input  io_rocc_dmem_0_acquire_valid,
    input [25:0] io_rocc_dmem_0_acquire_bits_addr_block,
    input [1:0] io_rocc_dmem_0_acquire_bits_client_xact_id,
    input [1:0] io_rocc_dmem_0_acquire_bits_addr_beat,
    input  io_rocc_dmem_0_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_dmem_0_acquire_bits_a_type,
    input [16:0] io_rocc_dmem_0_acquire_bits_union,
    input [127:0] io_rocc_dmem_0_acquire_bits_data,
    input  io_rocc_dmem_0_grant_ready,
    //output io_rocc_dmem_0_grant_valid
    //output[1:0] io_rocc_dmem_0_grant_bits_addr_beat
    //output[1:0] io_rocc_dmem_0_grant_bits_client_xact_id
    //output[3:0] io_rocc_dmem_0_grant_bits_manager_xact_id
    //output io_rocc_dmem_0_grant_bits_is_builtin_type
    //output[3:0] io_rocc_dmem_0_grant_bits_g_type
    //output[127:0] io_rocc_dmem_0_grant_bits_data
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [26:0] io_rocc_iptw_req_bits_addr,
    input [1:0] io_rocc_iptw_req_bits_prv,
    input  io_rocc_iptw_req_bits_store,
    input  io_rocc_iptw_req_bits_fetch,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[19:0] io_rocc_iptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_iptw_resp_bits_pte_reserved_for_software
    //output io_rocc_iptw_resp_bits_pte_d
    //output io_rocc_iptw_resp_bits_pte_r
    //output[3:0] io_rocc_iptw_resp_bits_pte_typ
    //output io_rocc_iptw_resp_bits_pte_v
    //output io_rocc_iptw_status_sd
    //output[30:0] io_rocc_iptw_status_zero2
    //output io_rocc_iptw_status_sd_rv32
    //output[8:0] io_rocc_iptw_status_zero1
    //output[4:0] io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_mprv
    //output[1:0] io_rocc_iptw_status_xs
    //output[1:0] io_rocc_iptw_status_fs
    //output[1:0] io_rocc_iptw_status_prv3
    //output io_rocc_iptw_status_ie3
    //output[1:0] io_rocc_iptw_status_prv2
    //output io_rocc_iptw_status_ie2
    //output[1:0] io_rocc_iptw_status_prv1
    //output io_rocc_iptw_status_ie1
    //output[1:0] io_rocc_iptw_status_prv
    //output io_rocc_iptw_status_ie
    //output io_rocc_iptw_invalidate
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [26:0] io_rocc_dptw_req_bits_addr,
    input [1:0] io_rocc_dptw_req_bits_prv,
    input  io_rocc_dptw_req_bits_store,
    input  io_rocc_dptw_req_bits_fetch,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[19:0] io_rocc_dptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_dptw_resp_bits_pte_reserved_for_software
    //output io_rocc_dptw_resp_bits_pte_d
    //output io_rocc_dptw_resp_bits_pte_r
    //output[3:0] io_rocc_dptw_resp_bits_pte_typ
    //output io_rocc_dptw_resp_bits_pte_v
    //output io_rocc_dptw_status_sd
    //output[30:0] io_rocc_dptw_status_zero2
    //output io_rocc_dptw_status_sd_rv32
    //output[8:0] io_rocc_dptw_status_zero1
    //output[4:0] io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_mprv
    //output[1:0] io_rocc_dptw_status_xs
    //output[1:0] io_rocc_dptw_status_fs
    //output[1:0] io_rocc_dptw_status_prv3
    //output io_rocc_dptw_status_ie3
    //output[1:0] io_rocc_dptw_status_prv2
    //output io_rocc_dptw_status_ie2
    //output[1:0] io_rocc_dptw_status_prv1
    //output io_rocc_dptw_status_ie1
    //output[1:0] io_rocc_dptw_status_prv
    //output io_rocc_dptw_status_ie
    //output io_rocc_dptw_invalidate
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [26:0] io_rocc_pptw_req_bits_addr,
    input [1:0] io_rocc_pptw_req_bits_prv,
    input  io_rocc_pptw_req_bits_store,
    input  io_rocc_pptw_req_bits_fetch,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[19:0] io_rocc_pptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_pptw_resp_bits_pte_reserved_for_software
    //output io_rocc_pptw_resp_bits_pte_d
    //output io_rocc_pptw_resp_bits_pte_r
    //output[3:0] io_rocc_pptw_resp_bits_pte_typ
    //output io_rocc_pptw_resp_bits_pte_v
    //output io_rocc_pptw_status_sd
    //output[30:0] io_rocc_pptw_status_zero2
    //output io_rocc_pptw_status_sd_rv32
    //output[8:0] io_rocc_pptw_status_zero1
    //output[4:0] io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_mprv
    //output[1:0] io_rocc_pptw_status_xs
    //output[1:0] io_rocc_pptw_status_fs
    //output[1:0] io_rocc_pptw_status_prv3
    //output io_rocc_pptw_status_ie3
    //output[1:0] io_rocc_pptw_status_prv2
    //output io_rocc_pptw_status_ie2
    //output[1:0] io_rocc_pptw_status_prv1
    //output io_rocc_pptw_status_ie1
    //output[1:0] io_rocc_pptw_status_prv
    //output io_rocc_pptw_status_ie
    //output io_rocc_pptw_invalidate
    //output io_rocc_exception
    output io_interrupt,
    output[63:0] io_interrupt_cause
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T882;
  wire csr_xcpt;
  wire insn_break;
  wire system_insn;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire insn_call;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire priv_sufficient;
  reg [1:0] reg_mstatus_prv;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  reg [1:0] reg_mstatus_prv1;
  wire[1:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  reg [1:0] reg_mstatus_prv2;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[63:0] wdata;
  wire[63:0] T38;
  wire[63:0] T39;
  reg [63:0] host_csr_bits_data;
  wire[63:0] T40;
  wire[63:0] T41;
  wire T42;
  wire host_csr_req_fire;
  wire T43;
  wire cpu_ren;
  wire T44;
  wire T45;
  reg  host_csr_req_valid;
  wire T46;
  wire T47;
  wire[63:0] T48;
  wire T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[11:0] addr;
  reg [11:0] host_csr_bits_addr;
  wire[11:0] T62;
  wire wen;
  wire T63;
  reg  host_csr_bits_rw;
  wire T64;
  wire T65;
  wire T66;
  wire read_only;
  wire[1:0] T67;
  wire cpu_wen;
  wire T68;
  wire T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[1:0] T883;
  wire T77;
  wire T78;
  wire T79;
  wire insn_ret;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire insn_redirect_trap;
  wire maybe_insn_redirect_trap;
  wire T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire[1:0] csr_addr_priv;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire fp_csr;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire addr_valid;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[2:0] T884;
  wire[3:0] T885;
  wire[1:0] T215;
  wire[1:0] T216;
  wire[1:0] T886;
  wire[63:0] T217;
  wire[63:0] T218;
  wire[63:0] T219;
  wire[63:0] T220;
  wire[63:0] T221;
  wire T222;
  wire T223;
  wire T224;
  reg  reg_mstatus_ie;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  reg  reg_mstatus_ie1;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  reg  reg_mstatus_ie2;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  reg  reg_mip_ssip;
  wire T887;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg  reg_mie_ssip;
  wire T888;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  reg  reg_mip_msip;
  wire T889;
  wire T265;
  wire T266;
  wire T267;
  reg  reg_mie_msip;
  wire T890;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  reg  reg_mip_stip;
  wire T891;
  wire T276;
  wire T277;
  reg  reg_mie_stip;
  wire T892;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  reg  reg_mip_mtip;
  wire T893;
  wire T288;
  wire T289;
  wire T290;
  reg [63:0] read_time;
  wire[63:0] T291;
  wire T292;
  reg [63:0] reg_mtimecmp;
  wire[63:0] T293;
  wire T294;
  reg  reg_mie_mtip;
  wire T894;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  reg [63:0] reg_fromhost;
  wire[63:0] T895;
  wire[63:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  reg [2:0] reg_frm;
  wire[2:0] T896;
  wire[63:0] T310;
  wire[63:0] T311;
  wire[63:0] T897;
  wire T312;
  wire[63:0] T898;
  wire[58:0] T313;
  wire T314;
  wire[63:0] T315;
  reg [5:0] R316;
  wire[5:0] T899;
  wire[5:0] T317;
  wire[6:0] T318;
  wire[6:0] T900;
  reg [57:0] R319;
  wire[57:0] T901;
  wire[57:0] T320;
  wire[57:0] T321;
  wire T322;
  wire insn_sfence_vm;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[39:0] T330;
  wire[39:0] T331;
  wire[39:0] T332;
  reg [39:0] reg_sepc;
  wire[39:0] T902;
  wire[63:0] T333;
  wire[63:0] T903;
  wire[39:0] T334;
  wire[63:0] T335;
  wire[63:0] T336;
  wire[63:0] T337;
  wire T338;
  reg [39:0] reg_mepc;
  wire[39:0] T904;
  wire[63:0] T339;
  wire[63:0] T905;
  wire[39:0] T340;
  wire[39:0] T341;
  wire[39:0] T342;
  wire[39:0] T343;
  wire[63:0] T344;
  wire[63:0] T345;
  wire[63:0] T346;
  wire T347;
  wire T348;
  wire[39:0] T349;
  reg [38:0] reg_stvec;
  wire[38:0] T906;
  wire[63:0] T350;
  wire[63:0] T907;
  wire[63:0] T351;
  wire[63:0] T352;
  wire[63:0] T353;
  wire T354;
  wire T355;
  wire[39:0] T908;
  wire[8:0] T356;
  wire[8:0] T909;
  wire[7:0] T357;
  wire T358;
  reg [31:0] reg_sptbr;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[19:0] T361;
  wire T362;
  reg  reg_mstatus_ie3;
  wire T363;
  reg [1:0] reg_mstatus_prv3;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[1:0] T910;
  wire T366;
  reg [1:0] reg_mstatus_fs;
  wire[1:0] T367;
  wire[1:0] T368;
  wire[1:0] T369;
  wire[1:0] T370;
  wire[1:0] T371;
  wire[1:0] T372;
  wire[1:0] T911;
  wire T373;
  reg [1:0] reg_mstatus_xs;
  wire[1:0] T374;
  reg  reg_mstatus_mprv;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  reg [4:0] reg_mstatus_vm;
  wire[4:0] T381;
  wire[4:0] T382;
  wire[4:0] T383;
  wire T384;
  wire T385;
  wire[4:0] T386;
  wire T387;
  wire T388;
  reg [8:0] reg_mstatus_zero1;
  wire[8:0] T389;
  reg  reg_mstatus_sd_rv32;
  wire T390;
  reg [30:0] reg_mstatus_zero2;
  wire[30:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  reg  reg_wfi;
  wire T912;
  wire T396;
  wire T397;
  wire insn_wfi;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire some_interrupt_pending;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire[63:0] T421;
  wire[63:0] T422;
  wire[63:0] T423;
  wire[24:0] T424;
  wire[24:0] T913;
  wire T425;
  wire[63:0] T426;
  wire[63:0] T427;
  wire[63:0] T428;
  wire[23:0] T429;
  wire[23:0] T914;
  wire T430;
  wire[63:0] T431;
  wire[63:0] T432;
  wire[63:0] T915;
  wire[31:0] T433;
  wire[63:0] T434;
  wire[63:0] T435;
  wire[63:0] T436;
  reg [39:0] reg_sbadaddr;
  wire[39:0] T437;
  reg [39:0] reg_mbadaddr;
  wire[39:0] T438;
  wire[39:0] T439;
  wire[39:0] T440;
  wire[39:0] T441;
  wire[38:0] T442;
  wire T443;
  wire T444;
  wire[24:0] T445;
  wire T446;
  wire T447;
  wire[38:0] T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire[39:0] T457;
  wire T458;
  wire[23:0] T459;
  wire[23:0] T916;
  wire T460;
  wire[63:0] T461;
  wire[63:0] T462;
  reg [63:0] reg_scause;
  wire[63:0] T463;
  reg [63:0] reg_mcause;
  wire[63:0] T464;
  wire[63:0] T465;
  wire[63:0] T466;
  wire[63:0] T467;
  wire[63:0] T468;
  wire T469;
  wire T470;
  wire[63:0] T917;
  wire[3:0] T471;
  wire[3:0] T918;
  wire T472;
  wire[63:0] T473;
  wire T474;
  wire[63:0] T475;
  wire[63:0] T476;
  reg [63:0] reg_sscratch;
  wire[63:0] T477;
  wire T478;
  wire[63:0] T479;
  wire[63:0] T919;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[3:0] T483;
  wire[1:0] T484;
  wire T485;
  wire T486;
  wire[1:0] T487;
  wire T488;
  wire T489;
  wire[3:0] T490;
  wire[1:0] T491;
  wire T492;
  wire T493;
  wire[1:0] T494;
  wire T495;
  wire T496;
  wire[63:0] T497;
  wire[63:0] T920;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[3:0] T501;
  wire[1:0] T502;
  wire T503;
  wire T504;
  wire[1:0] T505;
  wire T506;
  wire T507;
  wire[3:0] T508;
  wire[1:0] T509;
  wire T510;
  wire T511;
  wire[1:0] T512;
  wire T513;
  wire T514;
  wire[63:0] T515;
  wire[63:0] T516;
  wire[63:0] T517;
  wire[63:0] T518;
  wire[13:0] T519;
  wire[3:0] T520;
  wire[2:0] T521;
  wire T522;
  wire T523;
  wire[63:0] read_mstatus;
  wire[63:0] T524;
  wire[11:0] T525;
  wire[5:0] T526;
  wire[2:0] T527;
  wire[2:0] T528;
  wire[5:0] T529;
  wire[2:0] T530;
  wire[2:0] T531;
  wire[51:0] T532;
  wire[9:0] T533;
  wire[3:0] T534;
  wire[5:0] T535;
  wire[41:0] T536;
  wire[9:0] T537;
  wire[31:0] T538;
  wire[1:0] T539;
  wire T540;
  wire T541;
  wire[9:0] T542;
  wire[7:0] T543;
  wire T544;
  wire T545;
  wire[6:0] T546;
  wire[1:0] T547;
  wire[1:0] T548;
  wire[49:0] T549;
  wire[16:0] T550;
  wire[2:0] T551;
  wire[1:0] T552;
  wire[1:0] T553;
  wire T554;
  wire T555;
  wire[13:0] T556;
  wire[32:0] T557;
  wire[31:0] T558;
  wire T559;
  wire T560;
  wire[30:0] T561;
  wire T562;
  wire T563;
  wire[63:0] T564;
  wire[63:0] T565;
  wire[63:0] T566;
  reg [5:0] R567;
  wire[5:0] T921;
  wire[5:0] T568;
  wire[5:0] T569;
  wire[6:0] T570;
  wire[6:0] T922;
  wire T571;
  reg [57:0] R572;
  wire[57:0] T923;
  wire[57:0] T573;
  wire[57:0] T574;
  wire T575;
  wire T576;
  wire[63:0] T577;
  wire[63:0] T578;
  wire[63:0] T579;
  reg [5:0] R580;
  wire[5:0] T924;
  wire[5:0] T581;
  wire[5:0] T582;
  wire[6:0] T583;
  wire[6:0] T925;
  wire T584;
  reg [57:0] R585;
  wire[57:0] T926;
  wire[57:0] T586;
  wire[57:0] T587;
  wire T588;
  wire T589;
  wire[63:0] T590;
  wire[63:0] T591;
  wire[63:0] T592;
  reg [5:0] R593;
  wire[5:0] T927;
  wire[5:0] T594;
  wire[5:0] T595;
  wire[6:0] T596;
  wire[6:0] T928;
  wire T597;
  reg [57:0] R598;
  wire[57:0] T929;
  wire[57:0] T599;
  wire[57:0] T600;
  wire T601;
  wire T602;
  wire[63:0] T603;
  wire[63:0] T604;
  wire[63:0] T605;
  reg [5:0] R606;
  wire[5:0] T930;
  wire[5:0] T607;
  wire[5:0] T608;
  wire[6:0] T609;
  wire[6:0] T931;
  wire T610;
  reg [57:0] R611;
  wire[57:0] T932;
  wire[57:0] T612;
  wire[57:0] T613;
  wire T614;
  wire T615;
  wire[63:0] T616;
  wire[63:0] T617;
  wire[63:0] T618;
  reg [5:0] R619;
  wire[5:0] T933;
  wire[5:0] T620;
  wire[5:0] T621;
  wire[6:0] T622;
  wire[6:0] T934;
  wire T623;
  reg [57:0] R624;
  wire[57:0] T935;
  wire[57:0] T625;
  wire[57:0] T626;
  wire T627;
  wire T628;
  wire[63:0] T629;
  wire[63:0] T630;
  wire[63:0] T631;
  reg [5:0] R632;
  wire[5:0] T936;
  wire[5:0] T633;
  wire[5:0] T634;
  wire[6:0] T635;
  wire[6:0] T937;
  wire T636;
  reg [57:0] R637;
  wire[57:0] T938;
  wire[57:0] T638;
  wire[57:0] T639;
  wire T640;
  wire T641;
  wire[63:0] T642;
  wire[63:0] T643;
  wire[63:0] T644;
  reg [5:0] R645;
  wire[5:0] T939;
  wire[5:0] T646;
  wire[5:0] T647;
  wire[6:0] T648;
  wire[6:0] T940;
  wire T649;
  reg [57:0] R650;
  wire[57:0] T941;
  wire[57:0] T651;
  wire[57:0] T652;
  wire T653;
  wire T654;
  wire[63:0] T655;
  wire[63:0] T656;
  wire[63:0] T657;
  reg [5:0] R658;
  wire[5:0] T942;
  wire[5:0] T659;
  wire[5:0] T660;
  wire[6:0] T661;
  wire[6:0] T943;
  wire T662;
  reg [57:0] R663;
  wire[57:0] T944;
  wire[57:0] T664;
  wire[57:0] T665;
  wire T666;
  wire T667;
  wire[63:0] T668;
  wire[63:0] T669;
  wire[63:0] T670;
  reg [5:0] R671;
  wire[5:0] T945;
  wire[5:0] T672;
  wire[5:0] T673;
  wire[6:0] T674;
  wire[6:0] T946;
  wire T675;
  reg [57:0] R676;
  wire[57:0] T947;
  wire[57:0] T677;
  wire[57:0] T678;
  wire T679;
  wire T680;
  wire[63:0] T681;
  wire[63:0] T682;
  wire[63:0] T683;
  reg [5:0] R684;
  wire[5:0] T948;
  wire[5:0] T685;
  wire[5:0] T686;
  wire[6:0] T687;
  wire[6:0] T949;
  wire T688;
  reg [57:0] R689;
  wire[57:0] T950;
  wire[57:0] T690;
  wire[57:0] T691;
  wire T692;
  wire T693;
  wire[63:0] T694;
  wire[63:0] T695;
  wire[63:0] T696;
  reg [5:0] R697;
  wire[5:0] T951;
  wire[5:0] T698;
  wire[5:0] T699;
  wire[6:0] T700;
  wire[6:0] T952;
  wire T701;
  reg [57:0] R702;
  wire[57:0] T953;
  wire[57:0] T703;
  wire[57:0] T704;
  wire T705;
  wire T706;
  wire[63:0] T707;
  wire[63:0] T708;
  wire[63:0] T709;
  reg [5:0] R710;
  wire[5:0] T954;
  wire[5:0] T711;
  wire[5:0] T712;
  wire[6:0] T713;
  wire[6:0] T955;
  wire T714;
  reg [57:0] R715;
  wire[57:0] T956;
  wire[57:0] T716;
  wire[57:0] T717;
  wire T718;
  wire T719;
  wire[63:0] T720;
  wire[63:0] T721;
  wire[63:0] T722;
  reg [5:0] R723;
  wire[5:0] T957;
  wire[5:0] T724;
  wire[5:0] T725;
  wire[6:0] T726;
  wire[6:0] T958;
  wire T727;
  reg [57:0] R728;
  wire[57:0] T959;
  wire[57:0] T729;
  wire[57:0] T730;
  wire T731;
  wire T732;
  wire[63:0] T733;
  wire[63:0] T734;
  wire[63:0] T735;
  reg [5:0] R736;
  wire[5:0] T960;
  wire[5:0] T737;
  wire[5:0] T738;
  wire[6:0] T739;
  wire[6:0] T961;
  wire T740;
  reg [57:0] R741;
  wire[57:0] T962;
  wire[57:0] T742;
  wire[57:0] T743;
  wire T744;
  wire T745;
  wire[63:0] T746;
  wire[63:0] T747;
  wire[63:0] T748;
  reg [5:0] R749;
  wire[5:0] T963;
  wire[5:0] T750;
  wire[5:0] T751;
  wire[6:0] T752;
  wire[6:0] T964;
  wire T753;
  reg [57:0] R754;
  wire[57:0] T965;
  wire[57:0] T755;
  wire[57:0] T756;
  wire T757;
  wire T758;
  wire[63:0] T759;
  wire[63:0] T760;
  wire[63:0] T761;
  reg [5:0] R762;
  wire[5:0] T966;
  wire[5:0] T763;
  wire[5:0] T764;
  wire[6:0] T765;
  wire[6:0] T967;
  wire T766;
  reg [57:0] R767;
  wire[57:0] T968;
  wire[57:0] T768;
  wire[57:0] T769;
  wire T770;
  wire T771;
  wire[63:0] T772;
  wire[63:0] T773;
  wire[63:0] T774;
  reg [5:0] R775;
  wire[5:0] T969;
  wire[5:0] T776;
  wire[5:0] T777;
  wire[5:0] T778;
  wire[6:0] T779;
  wire[6:0] T970;
  wire T780;
  wire[5:0] T781;
  wire T782;
  reg [57:0] R783;
  wire[57:0] T971;
  wire[57:0] T784;
  wire[57:0] T785;
  wire[57:0] T786;
  wire T787;
  wire T788;
  wire[57:0] T789;
  wire[63:0] T790;
  wire[63:0] T791;
  wire[63:0] T792;
  wire[63:0] T793;
  wire[63:0] T794;
  wire[63:0] T795;
  reg [63:0] reg_tohost;
  wire[63:0] T972;
  wire[63:0] T796;
  wire[63:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire[63:0] T805;
  wire[63:0] T973;
  wire T806;
  reg  reg_stats;
  wire T974;
  wire T807;
  wire T808;
  wire T809;
  wire[63:0] T810;
  wire[63:0] T975;
  wire T811;
  wire[63:0] T812;
  wire[63:0] T976;
  wire T813;
  wire[63:0] T814;
  wire[63:0] T815;
  wire[63:0] T816;
  wire[63:0] T817;
  wire[63:0] T818;
  wire[63:0] T819;
  wire[63:0] T820;
  wire[23:0] T821;
  wire[23:0] T977;
  wire T822;
  wire[63:0] T823;
  wire[63:0] T824;
  wire[63:0] T825;
  wire[23:0] T826;
  wire[23:0] T978;
  wire T827;
  wire[63:0] T828;
  wire[63:0] T829;
  reg [63:0] reg_mscratch;
  wire[63:0] T830;
  wire T831;
  wire[63:0] T832;
  wire[63:0] T979;
  wire[7:0] T833;
  wire[7:0] T834;
  wire[7:0] T835;
  wire[3:0] T836;
  wire[1:0] T837;
  reg  reg_mie_usip;
  wire T980;
  wire[1:0] T838;
  reg  reg_mie_hsip;
  wire T981;
  wire[3:0] T839;
  wire[1:0] T840;
  reg  reg_mie_utip;
  wire T982;
  wire[1:0] T841;
  reg  reg_mie_htip;
  wire T983;
  wire[63:0] T842;
  wire[63:0] T984;
  wire[7:0] T843;
  wire[7:0] T844;
  wire[7:0] T845;
  wire[3:0] T846;
  wire[1:0] T847;
  reg  reg_mip_usip;
  wire T985;
  wire[1:0] T848;
  reg  reg_mip_hsip;
  wire T986;
  wire[3:0] T849;
  wire[1:0] T850;
  reg  reg_mip_utip;
  wire T987;
  wire[1:0] T851;
  reg  reg_mip_htip;
  wire T988;
  wire[63:0] T852;
  wire[63:0] T989;
  wire[8:0] T853;
  wire[63:0] T854;
  wire[63:0] T855;
  wire[63:0] T856;
  wire[63:0] T857;
  wire[63:0] T858;
  wire[63:0] T990;
  wire[63:0] T859;
  wire[63:0] T860;
  wire[63:0] T861;
  wire[63:0] T862;
  wire[63:0] T863;
  wire[63:0] T864;
  wire[63:0] T865;
  wire[63:0] T866;
  wire[63:0] T867;
  wire[63:0] T868;
  wire[63:0] T869;
  wire[63:0] T870;
  wire[63:0] T871;
  wire[63:0] T872;
  wire[63:0] T873;
  wire[63:0] T874;
  wire T991;
  wire T875;
  reg  host_csr_rep_valid;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    reg_mstatus_prv = {1{$random}};
    reg_mstatus_prv1 = {1{$random}};
    reg_mstatus_prv2 = {1{$random}};
    host_csr_bits_data = {2{$random}};
    host_csr_req_valid = {1{$random}};
    host_csr_bits_addr = {1{$random}};
    host_csr_bits_rw = {1{$random}};
    reg_mstatus_ie = {1{$random}};
    reg_mstatus_ie1 = {1{$random}};
    reg_mstatus_ie2 = {1{$random}};
    reg_mip_ssip = {1{$random}};
    reg_mie_ssip = {1{$random}};
    reg_mip_msip = {1{$random}};
    reg_mie_msip = {1{$random}};
    reg_mip_stip = {1{$random}};
    reg_mie_stip = {1{$random}};
    reg_mip_mtip = {1{$random}};
    read_time = {2{$random}};
    reg_mtimecmp = {2{$random}};
    reg_mie_mtip = {1{$random}};
    reg_fromhost = {2{$random}};
    reg_frm = {1{$random}};
    R316 = {1{$random}};
    R319 = {2{$random}};
    reg_sepc = {2{$random}};
    reg_mepc = {2{$random}};
    reg_stvec = {2{$random}};
    reg_sptbr = {1{$random}};
    reg_mstatus_ie3 = {1{$random}};
    reg_mstatus_prv3 = {1{$random}};
    reg_mstatus_fs = {1{$random}};
    reg_mstatus_xs = {1{$random}};
    reg_mstatus_mprv = {1{$random}};
    reg_mstatus_vm = {1{$random}};
    reg_mstatus_zero1 = {1{$random}};
    reg_mstatus_sd_rv32 = {1{$random}};
    reg_mstatus_zero2 = {1{$random}};
    reg_wfi = {1{$random}};
    reg_sbadaddr = {2{$random}};
    reg_mbadaddr = {2{$random}};
    reg_scause = {2{$random}};
    reg_mcause = {2{$random}};
    reg_sscratch = {2{$random}};
    R567 = {1{$random}};
    R572 = {2{$random}};
    R580 = {1{$random}};
    R585 = {2{$random}};
    R593 = {1{$random}};
    R598 = {2{$random}};
    R606 = {1{$random}};
    R611 = {2{$random}};
    R619 = {1{$random}};
    R624 = {2{$random}};
    R632 = {1{$random}};
    R637 = {2{$random}};
    R645 = {1{$random}};
    R650 = {2{$random}};
    R658 = {1{$random}};
    R663 = {2{$random}};
    R671 = {1{$random}};
    R676 = {2{$random}};
    R684 = {1{$random}};
    R689 = {2{$random}};
    R697 = {1{$random}};
    R702 = {2{$random}};
    R710 = {1{$random}};
    R715 = {2{$random}};
    R723 = {1{$random}};
    R728 = {2{$random}};
    R736 = {1{$random}};
    R741 = {2{$random}};
    R749 = {1{$random}};
    R754 = {2{$random}};
    R762 = {1{$random}};
    R767 = {2{$random}};
    R775 = {1{$random}};
    R783 = {2{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_mscratch = {2{$random}};
    reg_mie_usip = {1{$random}};
    reg_mie_hsip = {1{$random}};
    reg_mie_utip = {1{$random}};
    reg_mie_htip = {1{$random}};
    reg_mip_usip = {1{$random}};
    reg_mip_hsip = {1{$random}};
    reg_mip_utip = {1{$random}};
    reg_mip_htip = {1{$random}};
    host_csr_rep_valid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_rocc_exception = {1{$random}};
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_ie = {1{$random}};
//  assign io_rocc_pptw_status_prv = {1{$random}};
//  assign io_rocc_pptw_status_ie1 = {1{$random}};
//  assign io_rocc_pptw_status_prv1 = {1{$random}};
//  assign io_rocc_pptw_status_ie2 = {1{$random}};
//  assign io_rocc_pptw_status_prv2 = {1{$random}};
//  assign io_rocc_pptw_status_ie3 = {1{$random}};
//  assign io_rocc_pptw_status_prv3 = {1{$random}};
//  assign io_rocc_pptw_status_fs = {1{$random}};
//  assign io_rocc_pptw_status_xs = {1{$random}};
//  assign io_rocc_pptw_status_mprv = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_zero1 = {1{$random}};
//  assign io_rocc_pptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_pptw_status_zero2 = {1{$random}};
//  assign io_rocc_pptw_status_sd = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_ie = {1{$random}};
//  assign io_rocc_dptw_status_prv = {1{$random}};
//  assign io_rocc_dptw_status_ie1 = {1{$random}};
//  assign io_rocc_dptw_status_prv1 = {1{$random}};
//  assign io_rocc_dptw_status_ie2 = {1{$random}};
//  assign io_rocc_dptw_status_prv2 = {1{$random}};
//  assign io_rocc_dptw_status_ie3 = {1{$random}};
//  assign io_rocc_dptw_status_prv3 = {1{$random}};
//  assign io_rocc_dptw_status_fs = {1{$random}};
//  assign io_rocc_dptw_status_xs = {1{$random}};
//  assign io_rocc_dptw_status_mprv = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_zero1 = {1{$random}};
//  assign io_rocc_dptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_dptw_status_zero2 = {1{$random}};
//  assign io_rocc_dptw_status_sd = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_ie = {1{$random}};
//  assign io_rocc_iptw_status_prv = {1{$random}};
//  assign io_rocc_iptw_status_ie1 = {1{$random}};
//  assign io_rocc_iptw_status_prv1 = {1{$random}};
//  assign io_rocc_iptw_status_ie2 = {1{$random}};
//  assign io_rocc_iptw_status_prv2 = {1{$random}};
//  assign io_rocc_iptw_status_ie3 = {1{$random}};
//  assign io_rocc_iptw_status_prv3 = {1{$random}};
//  assign io_rocc_iptw_status_fs = {1{$random}};
//  assign io_rocc_iptw_status_xs = {1{$random}};
//  assign io_rocc_iptw_status_mprv = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_zero1 = {1{$random}};
//  assign io_rocc_iptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_iptw_status_zero2 = {1{$random}};
//  assign io_rocc_iptw_status_sd = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_data = {4{$random}};
//  assign io_rocc_dmem_0_grant_bits_g_type = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_dmem_0_grant_valid = {1{$random}};
//  assign io_rocc_dmem_0_acquire_ready = {1{$random}};
//  assign io_rocc_imem_grant_bits_data = {4{$random}};
//  assign io_rocc_imem_grant_bits_g_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_imem_grant_valid = {1{$random}};
//  assign io_rocc_imem_acquire_ready = {1{$random}};
//  assign io_rocc_s = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_data_word_bypass = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
//  assign io_rocc_cmd_bits_rs2 = {2{$random}};
//  assign io_rocc_cmd_bits_rs1 = {2{$random}};
//  assign io_rocc_cmd_bits_inst_opcode = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_funct = {1{$random}};
//  assign io_rocc_cmd_valid = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T3 <= 4'h1;
  assign T3 = T885 + T4;
  assign T4 = {1'h0, T5};
  assign T5 = T884 + T6;
  assign T6 = {1'h0, T7};
  assign T7 = T882 + T8;
  assign T8 = {1'h0, io_csr_replay};
  assign T882 = {1'h0, csr_xcpt};
  assign csr_xcpt = T13 | insn_break;
  assign insn_break = T9 & system_insn;
  assign system_insn = io_rw_cmd == 3'h4;
  assign T9 = T11 & T10;
  assign T10 = io_rw_addr[1'h0:1'h0];
  assign T11 = T12 ^ 1'h1;
  assign T12 = io_rw_addr[4'h8:4'h8];
  assign T13 = T19 | insn_call;
  assign insn_call = T14 & system_insn;
  assign T14 = T17 & T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = io_rw_addr[1'h0:1'h0];
  assign T17 = T18 ^ 1'h1;
  assign T18 = io_rw_addr[4'h8:4'h8];
  assign T19 = T96 | T20;
  assign T20 = system_insn & T21;
  assign T21 = priv_sufficient ^ 1'h1;
  assign priv_sufficient = csr_addr_priv <= reg_mstatus_prv;
  assign T22 = reset ? 2'h3 : T23;
  assign T23 = T90 ? T89 : T24;
  assign T24 = insn_redirect_trap ? 2'h1 : T25;
  assign T25 = insn_ret ? reg_mstatus_prv1 : T26;
  assign T26 = T27 ? 2'h3 : reg_mstatus_prv;
  assign T27 = io_exception | csr_xcpt;
  assign T28 = reset ? 2'h3 : T29;
  assign T29 = T78 ? T883 : T30;
  assign T30 = T71 ? T70 : T31;
  assign T31 = insn_ret ? reg_mstatus_prv2 : T32;
  assign T32 = T27 ? reg_mstatus_prv : reg_mstatus_prv1;
  assign T33 = reset ? 2'h0 : T34;
  assign T34 = T54 ? T37 : T35;
  assign T35 = insn_ret ? 2'h0 : T36;
  assign T36 = T27 ? reg_mstatus_prv1 : reg_mstatus_prv2;
  assign T37 = wdata[4'h8:3'h7];
  assign wdata = T53 ? io_rw_wdata : T38;
  assign T38 = T52 ? T50 : T39;
  assign T39 = T49 ? T48 : host_csr_bits_data;
  assign T40 = host_csr_req_fire ? io_rw_rdata : T41;
  assign T41 = T42 ? io_host_csr_req_bits_data : host_csr_bits_data;
  assign T42 = io_host_csr_req_ready & io_host_csr_req_valid;
  assign host_csr_req_fire = host_csr_req_valid & T43;
  assign T43 = cpu_ren ^ 1'h1;
  assign cpu_ren = T45 & T44;
  assign T44 = system_insn ^ 1'h1;
  assign T45 = io_rw_cmd != 3'h0;
  assign T46 = host_csr_req_fire ? 1'h0 : T47;
  assign T47 = T42 ? 1'h1 : host_csr_req_valid;
  assign T48 = io_rw_rdata | io_rw_wdata;
  assign T49 = io_rw_cmd == 3'h2;
  assign T50 = io_rw_rdata & T51;
  assign T51 = ~ io_rw_wdata;
  assign T52 = io_rw_cmd == 3'h3;
  assign T53 = io_rw_cmd == 3'h1;
  assign T54 = T60 & T55;
  assign T55 = T57 | T56;
  assign T56 = 2'h1 == T37;
  assign T57 = T59 | T58;
  assign T58 = 2'h0 == T37;
  assign T59 = 2'h3 == T37;
  assign T60 = wen & T61;
  assign T61 = addr == 12'h300;
  assign addr = cpu_ren ? io_rw_addr : host_csr_bits_addr;
  assign T62 = T42 ? io_host_csr_req_bits_addr : host_csr_bits_addr;
  assign wen = T65 | T63;
  assign T63 = host_csr_req_fire & host_csr_bits_rw;
  assign T64 = T42 ? io_host_csr_req_bits_rw : host_csr_bits_rw;
  assign T65 = cpu_wen & T66;
  assign T66 = read_only ^ 1'h1;
  assign read_only = T67 == 2'h3;
  assign T67 = io_rw_addr[4'hb:4'ha];
  assign cpu_wen = T68 & priv_sufficient;
  assign T68 = cpu_ren & T69;
  assign T69 = io_rw_cmd != 3'h5;
  assign T70 = wdata[3'h5:3'h4];
  assign T71 = T60 & T72;
  assign T72 = T74 | T73;
  assign T73 = 2'h1 == T70;
  assign T74 = T76 | T75;
  assign T75 = 2'h0 == T70;
  assign T76 = 2'h3 == T70;
  assign T883 = {1'h0, T77};
  assign T77 = wdata[3'h4:3'h4];
  assign T78 = wen & T79;
  assign T79 = addr == 12'h100;
  assign insn_ret = T80 & priv_sufficient;
  assign T80 = T81 & system_insn;
  assign T81 = T84 & T82;
  assign T82 = T83 ^ 1'h1;
  assign T83 = io_rw_addr[1'h0:1'h0];
  assign T84 = T87 & T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = io_rw_addr[1'h1:1'h1];
  assign T87 = io_rw_addr[4'h8:4'h8];
  assign insn_redirect_trap = maybe_insn_redirect_trap & priv_sufficient;
  assign maybe_insn_redirect_trap = T88 & system_insn;
  assign T88 = io_rw_addr[2'h2:2'h2];
  assign T89 = wdata[2'h2:1'h1];
  assign T90 = T60 & T91;
  assign T91 = T93 | T92;
  assign T92 = 2'h1 == T89;
  assign T93 = T95 | T94;
  assign T94 = 2'h0 == T89;
  assign T95 = 2'h3 == T89;
  assign csr_addr_priv = io_rw_addr[4'h9:4'h8];
  assign T96 = T214 | T97;
  assign T97 = cpu_ren & T98;
  assign T98 = T106 | T99;
  assign T99 = fp_csr & T100;
  assign T100 = T101 ^ 1'h1;
  assign T101 = io_status_fs != 2'h0;
  assign fp_csr = T103 | T102;
  assign T102 = addr == 12'h3;
  assign T103 = T105 | T104;
  assign T104 = addr == 12'h2;
  assign T105 = addr == 12'h1;
  assign T106 = T213 | T107;
  assign T107 = addr_valid ^ 1'h1;
  assign addr_valid = T109 | T108;
  assign T108 = addr == 12'h101;
  assign T109 = T111 | T110;
  assign T110 = addr == 12'h141;
  assign T111 = T113 | T112;
  assign T112 = addr == 12'h181;
  assign T113 = T115 | T114;
  assign T114 = addr == 12'h180;
  assign T115 = T117 | T116;
  assign T116 = addr == 12'hd43;
  assign T117 = T119 | T118;
  assign T118 = addr == 12'hd42;
  assign T119 = T121 | T120;
  assign T120 = addr == 12'h140;
  assign T121 = T123 | T122;
  assign T122 = addr == 12'h104;
  assign T123 = T125 | T124;
  assign T124 = addr == 12'h144;
  assign T125 = T126 | T79;
  assign T126 = T128 | T127;
  assign T127 = addr == 12'hccf;
  assign T128 = T130 | T129;
  assign T129 = addr == 12'hcce;
  assign T130 = T132 | T131;
  assign T131 = addr == 12'hccd;
  assign T132 = T134 | T133;
  assign T133 = addr == 12'hccc;
  assign T134 = T136 | T135;
  assign T135 = addr == 12'hccb;
  assign T136 = T138 | T137;
  assign T137 = addr == 12'hcca;
  assign T138 = T140 | T139;
  assign T139 = addr == 12'hcc9;
  assign T140 = T142 | T141;
  assign T141 = addr == 12'hcc8;
  assign T142 = T144 | T143;
  assign T143 = addr == 12'hcc7;
  assign T144 = T146 | T145;
  assign T145 = addr == 12'hcc6;
  assign T146 = T148 | T147;
  assign T147 = addr == 12'hcc5;
  assign T148 = T150 | T149;
  assign T149 = addr == 12'hcc4;
  assign T150 = T152 | T151;
  assign T151 = addr == 12'hcc3;
  assign T152 = T154 | T153;
  assign T153 = addr == 12'hcc2;
  assign T154 = T156 | T155;
  assign T155 = addr == 12'hcc1;
  assign T156 = T158 | T157;
  assign T157 = addr == 12'hcc0;
  assign T158 = T160 | T159;
  assign T159 = addr == 12'h902;
  assign T160 = T162 | T161;
  assign T161 = addr == 12'hc02;
  assign T162 = T164 | T163;
  assign T163 = addr == 12'h781;
  assign T164 = T166 | T165;
  assign T165 = addr == 12'h780;
  assign T166 = T168 | T167;
  assign T167 = addr == 12'hc0;
  assign T168 = T170 | T169;
  assign T169 = addr == 12'h783;
  assign T170 = T172 | T171;
  assign T171 = addr == 12'hf10;
  assign T172 = T174 | T173;
  assign T173 = addr == 12'h321;
  assign T174 = T176 | T175;
  assign T175 = addr == 12'h342;
  assign T176 = T178 | T177;
  assign T177 = addr == 12'h343;
  assign T178 = T180 | T179;
  assign T179 = addr == 12'h341;
  assign T180 = T182 | T181;
  assign T181 = addr == 12'h340;
  assign T182 = T184 | T183;
  assign T183 = addr == 12'h304;
  assign T184 = T186 | T185;
  assign T185 = addr == 12'h344;
  assign T186 = T188 | T187;
  assign T187 = addr == 12'h301;
  assign T188 = T190 | T189;
  assign T189 = addr == 12'h782;
  assign T190 = T192 | T191;
  assign T191 = addr == 12'h302;
  assign T192 = T193 | T61;
  assign T193 = T195 | T194;
  assign T194 = addr == 12'hf01;
  assign T195 = T197 | T196;
  assign T196 = addr == 12'hf00;
  assign T197 = T199 | T198;
  assign T198 = addr == 12'h701;
  assign T199 = T201 | T200;
  assign T200 = addr == 12'ha01;
  assign T201 = T203 | T202;
  assign T202 = addr == 12'hd01;
  assign T203 = T205 | T204;
  assign T204 = addr == 12'h901;
  assign T205 = T207 | T206;
  assign T206 = addr == 12'hc01;
  assign T207 = T209 | T208;
  assign T208 = addr == 12'h900;
  assign T209 = T211 | T210;
  assign T210 = addr == 12'hc00;
  assign T211 = T212 | T102;
  assign T212 = T105 | T104;
  assign T213 = priv_sufficient ^ 1'h1;
  assign T214 = cpu_wen & read_only;
  assign T884 = {2'h0, io_exception};
  assign T885 = {2'h0, T215};
  assign T215 = T886 + T216;
  assign T216 = {1'h0, insn_redirect_trap};
  assign T886 = {1'h0, insn_ret};
  assign io_interrupt_cause = T217;
  assign T217 = T297 ? 64'h8000000000000002 : T218;
  assign T218 = T282 ? 64'h8000000000000001 : T219;
  assign T219 = T270 ? 64'h8000000000000001 : T220;
  assign T220 = T259 ? 64'h8000000000000000 : T221;
  assign T221 = T222 ? 64'h8000000000000000 : 64'h0;
  assign T222 = T246 & T223;
  assign T223 = T245 | T224;
  assign T224 = T244 & reg_mstatus_ie;
  assign T225 = reset ? 1'h0 : T226;
  assign T226 = T78 ? T243 : T227;
  assign T227 = T60 ? T242 : T228;
  assign T228 = insn_ret ? reg_mstatus_ie1 : T229;
  assign T229 = T27 ? 1'h0 : reg_mstatus_ie;
  assign T230 = reset ? 1'h0 : T231;
  assign T231 = T78 ? T241 : T232;
  assign T232 = T60 ? T240 : T233;
  assign T233 = insn_ret ? reg_mstatus_ie2 : T234;
  assign T234 = T27 ? reg_mstatus_ie : reg_mstatus_ie1;
  assign T235 = reset ? 1'h0 : T236;
  assign T236 = T60 ? T239 : T237;
  assign T237 = insn_ret ? 1'h1 : T238;
  assign T238 = T27 ? reg_mstatus_ie1 : reg_mstatus_ie2;
  assign T239 = wdata[3'h6:3'h6];
  assign T240 = wdata[2'h3:2'h3];
  assign T241 = wdata[2'h3:2'h3];
  assign T242 = wdata[1'h0:1'h0];
  assign T243 = wdata[1'h0:1'h0];
  assign T244 = reg_mstatus_prv == 2'h1;
  assign T245 = reg_mstatus_prv < 2'h1;
  assign T246 = reg_mie_ssip & reg_mip_ssip;
  assign T887 = reset ? 1'h0 : T247;
  assign T247 = T252 ? T251 : T248;
  assign T248 = T250 ? T249 : reg_mip_ssip;
  assign T249 = wdata[1'h1:1'h1];
  assign T250 = wen & T185;
  assign T251 = wdata[1'h1:1'h1];
  assign T252 = wen & T124;
  assign T888 = reset ? 1'h0 : T253;
  assign T253 = T258 ? T257 : T254;
  assign T254 = T256 ? T255 : reg_mie_ssip;
  assign T255 = wdata[1'h1:1'h1];
  assign T256 = wen & T183;
  assign T257 = wdata[1'h1:1'h1];
  assign T258 = wen & T122;
  assign T259 = T264 & T260;
  assign T260 = T263 | T261;
  assign T261 = T262 & reg_mstatus_ie;
  assign T262 = reg_mstatus_prv == 2'h3;
  assign T263 = reg_mstatus_prv < 2'h3;
  assign T264 = reg_mie_msip & reg_mip_msip;
  assign T889 = reset ? 1'h0 : T265;
  assign T265 = io_host_ipi_rep_valid ? 1'h1 : T266;
  assign T266 = T250 ? T267 : reg_mip_msip;
  assign T267 = wdata[2'h3:2'h3];
  assign T890 = reset ? 1'h0 : T268;
  assign T268 = T256 ? T269 : reg_mie_msip;
  assign T269 = wdata[2'h3:2'h3];
  assign T270 = T275 & T271;
  assign T271 = T274 | T272;
  assign T272 = T273 & reg_mstatus_ie;
  assign T273 = reg_mstatus_prv == 2'h1;
  assign T274 = reg_mstatus_prv < 2'h1;
  assign T275 = reg_mie_stip & reg_mip_stip;
  assign T891 = reset ? 1'h0 : T276;
  assign T276 = T250 ? T277 : reg_mip_stip;
  assign T277 = wdata[3'h5:3'h5];
  assign T892 = reset ? 1'h0 : T278;
  assign T278 = T258 ? T281 : T279;
  assign T279 = T256 ? T280 : reg_mie_stip;
  assign T280 = wdata[3'h5:3'h5];
  assign T281 = wdata[3'h5:3'h5];
  assign T282 = T287 & T283;
  assign T283 = T286 | T284;
  assign T284 = T285 & reg_mstatus_ie;
  assign T285 = reg_mstatus_prv == 2'h3;
  assign T286 = reg_mstatus_prv < 2'h3;
  assign T287 = reg_mie_mtip & reg_mip_mtip;
  assign T893 = reset ? 1'h0 : T288;
  assign T288 = T294 ? 1'h0 : T289;
  assign T289 = T290 ? 1'h1 : reg_mip_mtip;
  assign T290 = reg_mtimecmp <= read_time;
  assign T291 = T292 ? wdata : read_time;
  assign T292 = wen & T198;
  assign T293 = T294 ? wdata : reg_mtimecmp;
  assign T294 = wen & T173;
  assign T894 = reset ? 1'h0 : T295;
  assign T295 = T256 ? T296 : reg_mie_mtip;
  assign T296 = wdata[3'h7:3'h7];
  assign T297 = T302 & T298;
  assign T298 = T301 | T299;
  assign T299 = T300 & reg_mstatus_ie;
  assign T300 = reg_mstatus_prv == 2'h3;
  assign T301 = reg_mstatus_prv < 2'h3;
  assign T302 = reg_fromhost != 64'h0;
  assign T895 = reset ? 64'h0 : T303;
  assign T303 = T304 ? wdata : reg_fromhost;
  assign T304 = T308 & T305;
  assign T305 = T307 | T306;
  assign T306 = host_csr_req_fire ^ 1'h1;
  assign T307 = reg_fromhost == 64'h0;
  assign T308 = wen & T163;
  assign io_interrupt = T309;
  assign T309 = io_interrupt_cause[6'h3f:6'h3f];
  assign io_fcsr_rm = reg_frm;
  assign T896 = T310[2'h2:1'h0];
  assign T310 = T314 ? T898 : T311;
  assign T311 = T312 ? wdata : T897;
  assign T897 = {61'h0, reg_frm};
  assign T312 = wen & T104;
  assign T898 = {5'h0, T313};
  assign T313 = wdata >> 3'h5;
  assign T314 = wen & T102;
  assign io_time = T315;
  assign T315 = {R319, R316};
  assign T899 = reset ? 6'h0 : T317;
  assign T317 = T318[3'h5:1'h0];
  assign T318 = T900 + 7'h1;
  assign T900 = {1'h0, R316};
  assign T901 = reset ? 58'h0 : T320;
  assign T320 = T322 ? T321 : R319;
  assign T321 = R319 + 58'h1;
  assign T322 = T318[3'h6:3'h6];
  assign io_fatc = insn_sfence_vm;
  assign insn_sfence_vm = T323 & priv_sufficient;
  assign T323 = T324 & system_insn;
  assign T324 = T326 & T325;
  assign T325 = io_rw_addr[1'h0:1'h0];
  assign T326 = T329 & T327;
  assign T327 = T328 ^ 1'h1;
  assign T328 = io_rw_addr[1'h1:1'h1];
  assign T329 = io_rw_addr[4'h8:4'h8];
  assign io_evec = T330;
  assign T330 = T358 ? T908 : T331;
  assign T331 = maybe_insn_redirect_trap ? T349 : T332;
  assign T332 = T348 ? reg_mepc : reg_sepc;
  assign T902 = T333[6'h27:1'h0];
  assign T333 = T338 ? T335 : T903;
  assign T903 = {24'h0, T334};
  assign T334 = insn_redirect_trap ? reg_mepc : reg_sepc;
  assign T335 = ~ T336;
  assign T336 = T337 | 64'h3;
  assign T337 = ~ wdata;
  assign T338 = wen & T110;
  assign T904 = T339[6'h27:1'h0];
  assign T339 = T347 ? T344 : T905;
  assign T905 = {24'h0, T340};
  assign T340 = T27 ? T341 : reg_mepc;
  assign T341 = ~ T342;
  assign T342 = T343 | 40'h3;
  assign T343 = ~ io_pc;
  assign T344 = ~ T345;
  assign T345 = T346 | 64'h3;
  assign T346 = ~ wdata;
  assign T347 = wen & T179;
  assign T348 = reg_mstatus_prv[1'h1:1'h1];
  assign T349 = {T355, reg_stvec};
  assign T906 = T350[6'h26:1'h0];
  assign T350 = T354 ? T351 : T907;
  assign T907 = {25'h0, reg_stvec};
  assign T351 = ~ T352;
  assign T352 = T353 | 64'h3;
  assign T353 = ~ wdata;
  assign T354 = wen & T108;
  assign T355 = reg_stvec[6'h26:6'h26];
  assign T908 = {31'h0, T356};
  assign T356 = T909 + 9'h100;
  assign T909 = {1'h0, T357};
  assign T357 = reg_mstatus_prv << 3'h6;
  assign T358 = io_exception | csr_xcpt;
  assign io_ptbr = reg_sptbr;
  assign T359 = T362 ? T360 : reg_sptbr;
  assign T360 = {T361, 12'h0};
  assign T361 = wdata[5'h1f:4'hc];
  assign T362 = wen & T114;
  assign io_status_ie = reg_mstatus_ie;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_ie1 = reg_mstatus_ie1;
  assign io_status_prv1 = reg_mstatus_prv1;
  assign io_status_ie2 = reg_mstatus_ie2;
  assign io_status_prv2 = reg_mstatus_prv2;
  assign io_status_ie3 = reg_mstatus_ie3;
  assign T363 = reset ? 1'h0 : reg_mstatus_ie3;
  assign io_status_prv3 = reg_mstatus_prv3;
  assign T364 = reset ? 2'h0 : reg_mstatus_prv3;
  assign io_status_fs = T365;
  assign T365 = 2'h0 - T910;
  assign T910 = {1'h0, T366};
  assign T366 = reg_mstatus_fs != 2'h0;
  assign T367 = reset ? 2'h0 : T368;
  assign T368 = T78 ? T371 : T369;
  assign T369 = T60 ? T370 : reg_mstatus_fs;
  assign T370 = wdata[4'hd:4'hc];
  assign T371 = wdata[4'hd:4'hc];
  assign io_status_xs = T372;
  assign T372 = 2'h0 - T911;
  assign T911 = {1'h0, T373};
  assign T373 = reg_mstatus_xs != 2'h0;
  assign T374 = reset ? 2'h0 : reg_mstatus_xs;
  assign io_status_mprv = reg_mstatus_mprv;
  assign T375 = reset ? 1'h0 : T376;
  assign T376 = T78 ? T380 : T377;
  assign T377 = T60 ? T379 : T378;
  assign T378 = T27 ? 1'h0 : reg_mstatus_mprv;
  assign T379 = wdata[5'h10:5'h10];
  assign T380 = wdata[5'h10:5'h10];
  assign io_status_vm = reg_mstatus_vm;
  assign T381 = reset ? 5'h0 : T382;
  assign T382 = T387 ? 5'h9 : T383;
  assign T383 = T384 ? 5'h0 : reg_mstatus_vm;
  assign T384 = T60 & T385;
  assign T385 = T386 == 5'h0;
  assign T386 = wdata[5'h15:5'h11];
  assign T387 = T60 & T388;
  assign T388 = T386 == 5'h9;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign T389 = reset ? 9'h0 : reg_mstatus_zero1;
  assign io_status_sd_rv32 = reg_mstatus_sd_rv32;
  assign T390 = reset ? 1'h0 : reg_mstatus_sd_rv32;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign T391 = reset ? 31'h0 : reg_mstatus_zero2;
  assign io_status_sd = T392;
  assign T392 = T394 | T393;
  assign T393 = io_status_xs == 2'h3;
  assign T394 = io_status_fs == 2'h3;
  assign io_eret = T395;
  assign T395 = insn_ret | insn_redirect_trap;
  assign io_csr_xcpt = csr_xcpt;
  assign io_csr_stall = reg_wfi;
  assign T912 = reset ? 1'h0 : T396;
  assign T396 = some_interrupt_pending ? 1'h0 : T397;
  assign T397 = insn_wfi ? 1'h1 : reg_wfi;
  assign insn_wfi = T398 & priv_sufficient;
  assign T398 = T399 & system_insn;
  assign T399 = T402 & T400;
  assign T400 = T401 ^ 1'h1;
  assign T401 = io_rw_addr[1'h0:1'h0];
  assign T402 = T404 & T403;
  assign T403 = io_rw_addr[1'h1:1'h1];
  assign T404 = io_rw_addr[4'h8:4'h8];
  assign some_interrupt_pending = T405;
  assign T405 = T417 ? 1'h1 : T406;
  assign T406 = T415 ? 1'h1 : T407;
  assign T407 = T413 ? 1'h1 : T408;
  assign T408 = T411 ? 1'h1 : T409;
  assign T409 = T246 & T410;
  assign T410 = reg_mstatus_prv <= 2'h1;
  assign T411 = T264 & T412;
  assign T412 = reg_mstatus_prv <= 2'h3;
  assign T413 = T275 & T414;
  assign T414 = reg_mstatus_prv <= 2'h1;
  assign T415 = T287 & T416;
  assign T416 = reg_mstatus_prv <= 2'h3;
  assign T417 = T302 & T418;
  assign T418 = reg_mstatus_prv <= 2'h3;
  assign io_csr_replay = T419;
  assign T419 = io_host_ipi_req_valid & T420;
  assign T420 = io_host_ipi_req_ready ^ 1'h1;
  assign io_rw_rdata = T421;
  assign T421 = T426 | T422;
  assign T422 = T108 ? T423 : 64'h0;
  assign T423 = {T424, reg_stvec};
  assign T424 = 25'h0 - T913;
  assign T913 = {24'h0, T425};
  assign T425 = reg_stvec[6'h26:6'h26];
  assign T426 = T431 | T427;
  assign T427 = T110 ? T428 : 64'h0;
  assign T428 = {T429, reg_sepc};
  assign T429 = 24'h0 - T914;
  assign T914 = {23'h0, T430};
  assign T430 = reg_sepc[6'h27:6'h27];
  assign T431 = T432 | 64'h0;
  assign T432 = T434 | T915;
  assign T915 = {32'h0, T433};
  assign T433 = T114 ? reg_sptbr : 32'h0;
  assign T434 = T461 | T435;
  assign T435 = T116 ? T436 : 64'h0;
  assign T436 = {T459, reg_sbadaddr};
  assign T437 = insn_redirect_trap ? reg_mbadaddr : reg_sbadaddr;
  assign T438 = T458 ? T457 : T439;
  assign T439 = T449 ? T441 : T440;
  assign T440 = T27 ? io_pc : reg_mbadaddr;
  assign T441 = {T443, T442};
  assign T442 = io_rw_wdata[6'h26:1'h0];
  assign T443 = T447 ? T446 : T444;
  assign T444 = T445 != 25'h0;
  assign T445 = io_rw_wdata[6'h3f:6'h27];
  assign T446 = T445 == 25'h1ffffff;
  assign T447 = $signed(T448) < $signed(1'h0);
  assign T448 = T442;
  assign T449 = T27 & T450;
  assign T450 = T452 | T451;
  assign T451 = io_cause == 64'h6;
  assign T452 = T454 | T453;
  assign T453 = io_cause == 64'h7;
  assign T454 = T456 | T455;
  assign T455 = io_cause == 64'h4;
  assign T456 = io_cause == 64'h5;
  assign T457 = wdata[6'h27:1'h0];
  assign T458 = wen & T177;
  assign T459 = 24'h0 - T916;
  assign T916 = {23'h0, T460};
  assign T460 = reg_sbadaddr[6'h27:6'h27];
  assign T461 = T475 | T462;
  assign T462 = T118 ? reg_scause : 64'h0;
  assign T463 = insn_redirect_trap ? reg_mcause : reg_scause;
  assign T464 = T474 ? T473 : T465;
  assign T465 = T472 ? T917 : T466;
  assign T466 = T470 ? 64'h3 : T467;
  assign T467 = T469 ? 64'h2 : T468;
  assign T468 = T27 ? io_cause : reg_mcause;
  assign T469 = T27 & csr_xcpt;
  assign T470 = T469 & insn_break;
  assign T917 = {60'h0, T471};
  assign T471 = T918 + 4'h8;
  assign T918 = {2'h0, reg_mstatus_prv};
  assign T472 = T469 & insn_call;
  assign T473 = wdata & 64'h800000000000001f;
  assign T474 = wen & T175;
  assign T475 = T479 | T476;
  assign T476 = T120 ? reg_sscratch : 64'h0;
  assign T477 = T478 ? wdata : reg_sscratch;
  assign T478 = wen & T120;
  assign T479 = T497 | T919;
  assign T919 = {56'h0, T480};
  assign T480 = T122 ? T481 : 8'h0;
  assign T481 = T482;
  assign T482 = {T490, T483};
  assign T483 = {T487, T484};
  assign T484 = {T486, T485};
  assign T485 = 1'h0;
  assign T486 = reg_mie_ssip;
  assign T487 = {T489, T488};
  assign T488 = 1'h0;
  assign T489 = 1'h0;
  assign T490 = {T494, T491};
  assign T491 = {T493, T492};
  assign T492 = 1'h0;
  assign T493 = reg_mie_stip;
  assign T494 = {T496, T495};
  assign T495 = 1'h0;
  assign T496 = 1'h0;
  assign T497 = T515 | T920;
  assign T920 = {56'h0, T498};
  assign T498 = T124 ? T499 : 8'h0;
  assign T499 = T500;
  assign T500 = {T508, T501};
  assign T501 = {T505, T502};
  assign T502 = {T504, T503};
  assign T503 = 1'h0;
  assign T504 = reg_mip_ssip;
  assign T505 = {T507, T506};
  assign T506 = 1'h0;
  assign T507 = 1'h0;
  assign T508 = {T512, T509};
  assign T509 = {T511, T510};
  assign T510 = 1'h0;
  assign T511 = reg_mip_stip;
  assign T512 = {T514, T513};
  assign T513 = 1'h0;
  assign T514 = 1'h0;
  assign T515 = T564 | T516;
  assign T516 = T79 ? T517 : 64'h0;
  assign T517 = T518;
  assign T518 = {T549, T519};
  assign T519 = {T542, T520};
  assign T520 = {T540, T521};
  assign T521 = {T539, T522};
  assign T522 = T523;
  assign T523 = read_mstatus[1'h0:1'h0];
  assign read_mstatus = T524;
  assign T524 = {T532, T525};
  assign T525 = {T529, T526};
  assign T526 = {T528, T527};
  assign T527 = {io_status_prv, io_status_ie};
  assign T528 = {io_status_prv1, io_status_ie1};
  assign T529 = {T531, T530};
  assign T530 = {io_status_prv2, io_status_ie2};
  assign T531 = {io_status_prv3, io_status_ie3};
  assign T532 = {T536, T533};
  assign T533 = {T535, T534};
  assign T534 = {io_status_xs, io_status_fs};
  assign T535 = {io_status_vm, io_status_mprv};
  assign T536 = {T538, T537};
  assign T537 = {io_status_sd_rv32, io_status_zero1};
  assign T538 = {io_status_sd, io_status_zero2};
  assign T539 = 2'h0;
  assign T540 = T541;
  assign T541 = read_mstatus[2'h3:2'h3];
  assign T542 = {T547, T543};
  assign T543 = {T546, T544};
  assign T544 = T545;
  assign T545 = read_mstatus[3'h4:3'h4];
  assign T546 = 7'h0;
  assign T547 = T548;
  assign T548 = read_mstatus[4'hd:4'hc];
  assign T549 = {T557, T550};
  assign T550 = {T556, T551};
  assign T551 = {T554, T552};
  assign T552 = T553;
  assign T553 = read_mstatus[4'hf:4'he];
  assign T554 = T555;
  assign T555 = read_mstatus[5'h10:5'h10];
  assign T556 = 14'h0;
  assign T557 = {T562, T558};
  assign T558 = {T561, T559};
  assign T559 = T560;
  assign T560 = read_mstatus[5'h1f:5'h1f];
  assign T561 = 31'h0;
  assign T562 = T563;
  assign T563 = read_mstatus[6'h3f:6'h3f];
  assign T564 = T577 | T565;
  assign T565 = T127 ? T566 : 64'h0;
  assign T566 = {R572, R567};
  assign T921 = reset ? 6'h0 : T568;
  assign T568 = T571 ? T569 : R567;
  assign T569 = T570[3'h5:1'h0];
  assign T570 = T922 + 7'h1;
  assign T922 = {1'h0, R567};
  assign T571 = io_uarch_counters_15 != 1'h0;
  assign T923 = reset ? 58'h0 : T573;
  assign T573 = T575 ? T574 : R572;
  assign T574 = R572 + 58'h1;
  assign T575 = T571 & T576;
  assign T576 = T570[3'h6:3'h6];
  assign T577 = T590 | T578;
  assign T578 = T129 ? T579 : 64'h0;
  assign T579 = {R585, R580};
  assign T924 = reset ? 6'h0 : T581;
  assign T581 = T584 ? T582 : R580;
  assign T582 = T583[3'h5:1'h0];
  assign T583 = T925 + 7'h1;
  assign T925 = {1'h0, R580};
  assign T584 = io_uarch_counters_14 != 1'h0;
  assign T926 = reset ? 58'h0 : T586;
  assign T586 = T588 ? T587 : R585;
  assign T587 = R585 + 58'h1;
  assign T588 = T584 & T589;
  assign T589 = T583[3'h6:3'h6];
  assign T590 = T603 | T591;
  assign T591 = T131 ? T592 : 64'h0;
  assign T592 = {R598, R593};
  assign T927 = reset ? 6'h0 : T594;
  assign T594 = T597 ? T595 : R593;
  assign T595 = T596[3'h5:1'h0];
  assign T596 = T928 + 7'h1;
  assign T928 = {1'h0, R593};
  assign T597 = io_uarch_counters_13 != 1'h0;
  assign T929 = reset ? 58'h0 : T599;
  assign T599 = T601 ? T600 : R598;
  assign T600 = R598 + 58'h1;
  assign T601 = T597 & T602;
  assign T602 = T596[3'h6:3'h6];
  assign T603 = T616 | T604;
  assign T604 = T133 ? T605 : 64'h0;
  assign T605 = {R611, R606};
  assign T930 = reset ? 6'h0 : T607;
  assign T607 = T610 ? T608 : R606;
  assign T608 = T609[3'h5:1'h0];
  assign T609 = T931 + 7'h1;
  assign T931 = {1'h0, R606};
  assign T610 = io_uarch_counters_12 != 1'h0;
  assign T932 = reset ? 58'h0 : T612;
  assign T612 = T614 ? T613 : R611;
  assign T613 = R611 + 58'h1;
  assign T614 = T610 & T615;
  assign T615 = T609[3'h6:3'h6];
  assign T616 = T629 | T617;
  assign T617 = T135 ? T618 : 64'h0;
  assign T618 = {R624, R619};
  assign T933 = reset ? 6'h0 : T620;
  assign T620 = T623 ? T621 : R619;
  assign T621 = T622[3'h5:1'h0];
  assign T622 = T934 + 7'h1;
  assign T934 = {1'h0, R619};
  assign T623 = io_uarch_counters_11 != 1'h0;
  assign T935 = reset ? 58'h0 : T625;
  assign T625 = T627 ? T626 : R624;
  assign T626 = R624 + 58'h1;
  assign T627 = T623 & T628;
  assign T628 = T622[3'h6:3'h6];
  assign T629 = T642 | T630;
  assign T630 = T137 ? T631 : 64'h0;
  assign T631 = {R637, R632};
  assign T936 = reset ? 6'h0 : T633;
  assign T633 = T636 ? T634 : R632;
  assign T634 = T635[3'h5:1'h0];
  assign T635 = T937 + 7'h1;
  assign T937 = {1'h0, R632};
  assign T636 = io_uarch_counters_10 != 1'h0;
  assign T938 = reset ? 58'h0 : T638;
  assign T638 = T640 ? T639 : R637;
  assign T639 = R637 + 58'h1;
  assign T640 = T636 & T641;
  assign T641 = T635[3'h6:3'h6];
  assign T642 = T655 | T643;
  assign T643 = T139 ? T644 : 64'h0;
  assign T644 = {R650, R645};
  assign T939 = reset ? 6'h0 : T646;
  assign T646 = T649 ? T647 : R645;
  assign T647 = T648[3'h5:1'h0];
  assign T648 = T940 + 7'h1;
  assign T940 = {1'h0, R645};
  assign T649 = io_uarch_counters_9 != 1'h0;
  assign T941 = reset ? 58'h0 : T651;
  assign T651 = T653 ? T652 : R650;
  assign T652 = R650 + 58'h1;
  assign T653 = T649 & T654;
  assign T654 = T648[3'h6:3'h6];
  assign T655 = T668 | T656;
  assign T656 = T141 ? T657 : 64'h0;
  assign T657 = {R663, R658};
  assign T942 = reset ? 6'h0 : T659;
  assign T659 = T662 ? T660 : R658;
  assign T660 = T661[3'h5:1'h0];
  assign T661 = T943 + 7'h1;
  assign T943 = {1'h0, R658};
  assign T662 = io_uarch_counters_8 != 1'h0;
  assign T944 = reset ? 58'h0 : T664;
  assign T664 = T666 ? T665 : R663;
  assign T665 = R663 + 58'h1;
  assign T666 = T662 & T667;
  assign T667 = T661[3'h6:3'h6];
  assign T668 = T681 | T669;
  assign T669 = T143 ? T670 : 64'h0;
  assign T670 = {R676, R671};
  assign T945 = reset ? 6'h0 : T672;
  assign T672 = T675 ? T673 : R671;
  assign T673 = T674[3'h5:1'h0];
  assign T674 = T946 + 7'h1;
  assign T946 = {1'h0, R671};
  assign T675 = io_uarch_counters_7 != 1'h0;
  assign T947 = reset ? 58'h0 : T677;
  assign T677 = T679 ? T678 : R676;
  assign T678 = R676 + 58'h1;
  assign T679 = T675 & T680;
  assign T680 = T674[3'h6:3'h6];
  assign T681 = T694 | T682;
  assign T682 = T145 ? T683 : 64'h0;
  assign T683 = {R689, R684};
  assign T948 = reset ? 6'h0 : T685;
  assign T685 = T688 ? T686 : R684;
  assign T686 = T687[3'h5:1'h0];
  assign T687 = T949 + 7'h1;
  assign T949 = {1'h0, R684};
  assign T688 = io_uarch_counters_6 != 1'h0;
  assign T950 = reset ? 58'h0 : T690;
  assign T690 = T692 ? T691 : R689;
  assign T691 = R689 + 58'h1;
  assign T692 = T688 & T693;
  assign T693 = T687[3'h6:3'h6];
  assign T694 = T707 | T695;
  assign T695 = T147 ? T696 : 64'h0;
  assign T696 = {R702, R697};
  assign T951 = reset ? 6'h0 : T698;
  assign T698 = T701 ? T699 : R697;
  assign T699 = T700[3'h5:1'h0];
  assign T700 = T952 + 7'h1;
  assign T952 = {1'h0, R697};
  assign T701 = io_uarch_counters_5 != 1'h0;
  assign T953 = reset ? 58'h0 : T703;
  assign T703 = T705 ? T704 : R702;
  assign T704 = R702 + 58'h1;
  assign T705 = T701 & T706;
  assign T706 = T700[3'h6:3'h6];
  assign T707 = T720 | T708;
  assign T708 = T149 ? T709 : 64'h0;
  assign T709 = {R715, R710};
  assign T954 = reset ? 6'h0 : T711;
  assign T711 = T714 ? T712 : R710;
  assign T712 = T713[3'h5:1'h0];
  assign T713 = T955 + 7'h1;
  assign T955 = {1'h0, R710};
  assign T714 = io_uarch_counters_4 != 1'h0;
  assign T956 = reset ? 58'h0 : T716;
  assign T716 = T718 ? T717 : R715;
  assign T717 = R715 + 58'h1;
  assign T718 = T714 & T719;
  assign T719 = T713[3'h6:3'h6];
  assign T720 = T733 | T721;
  assign T721 = T151 ? T722 : 64'h0;
  assign T722 = {R728, R723};
  assign T957 = reset ? 6'h0 : T724;
  assign T724 = T727 ? T725 : R723;
  assign T725 = T726[3'h5:1'h0];
  assign T726 = T958 + 7'h1;
  assign T958 = {1'h0, R723};
  assign T727 = io_uarch_counters_3 != 1'h0;
  assign T959 = reset ? 58'h0 : T729;
  assign T729 = T731 ? T730 : R728;
  assign T730 = R728 + 58'h1;
  assign T731 = T727 & T732;
  assign T732 = T726[3'h6:3'h6];
  assign T733 = T746 | T734;
  assign T734 = T153 ? T735 : 64'h0;
  assign T735 = {R741, R736};
  assign T960 = reset ? 6'h0 : T737;
  assign T737 = T740 ? T738 : R736;
  assign T738 = T739[3'h5:1'h0];
  assign T739 = T961 + 7'h1;
  assign T961 = {1'h0, R736};
  assign T740 = io_uarch_counters_2 != 1'h0;
  assign T962 = reset ? 58'h0 : T742;
  assign T742 = T744 ? T743 : R741;
  assign T743 = R741 + 58'h1;
  assign T744 = T740 & T745;
  assign T745 = T739[3'h6:3'h6];
  assign T746 = T759 | T747;
  assign T747 = T155 ? T748 : 64'h0;
  assign T748 = {R754, R749};
  assign T963 = reset ? 6'h0 : T750;
  assign T750 = T753 ? T751 : R749;
  assign T751 = T752[3'h5:1'h0];
  assign T752 = T964 + 7'h1;
  assign T964 = {1'h0, R749};
  assign T753 = io_uarch_counters_1 != 1'h0;
  assign T965 = reset ? 58'h0 : T755;
  assign T755 = T757 ? T756 : R754;
  assign T756 = R754 + 58'h1;
  assign T757 = T753 & T758;
  assign T758 = T752[3'h6:3'h6];
  assign T759 = T772 | T760;
  assign T760 = T157 ? T761 : 64'h0;
  assign T761 = {R767, R762};
  assign T966 = reset ? 6'h0 : T763;
  assign T763 = T766 ? T764 : R762;
  assign T764 = T765[3'h5:1'h0];
  assign T765 = T967 + 7'h1;
  assign T967 = {1'h0, R762};
  assign T766 = io_uarch_counters_0 != 1'h0;
  assign T968 = reset ? 58'h0 : T768;
  assign T768 = T770 ? T769 : R767;
  assign T769 = R767 + 58'h1;
  assign T770 = T766 & T771;
  assign T771 = T765[3'h6:3'h6];
  assign T772 = T790 | T773;
  assign T773 = T159 ? T774 : 64'h0;
  assign T774 = {R783, R775};
  assign T969 = reset ? 6'h0 : T776;
  assign T776 = T782 ? T781 : T777;
  assign T777 = T780 ? T778 : R775;
  assign T778 = T779[3'h5:1'h0];
  assign T779 = T970 + 7'h1;
  assign T970 = {1'h0, R775};
  assign T780 = io_retire != 1'h0;
  assign T781 = wdata[3'h5:1'h0];
  assign T782 = wen & T159;
  assign T971 = reset ? 58'h0 : T784;
  assign T784 = T782 ? T789 : T785;
  assign T785 = T787 ? T786 : R783;
  assign T786 = R783 + 58'h1;
  assign T787 = T780 & T788;
  assign T788 = T779[3'h6:3'h6];
  assign T789 = wdata[6'h3f:3'h6];
  assign T790 = T792 | T791;
  assign T791 = T161 ? T774 : 64'h0;
  assign T792 = T794 | T793;
  assign T793 = T163 ? reg_fromhost : 64'h0;
  assign T794 = T805 | T795;
  assign T795 = T165 ? reg_tohost : 64'h0;
  assign T972 = reset ? 64'h0 : T796;
  assign T796 = T801 ? wdata : T797;
  assign T797 = T798 ? 64'h0 : reg_tohost;
  assign T798 = T799 & T165;
  assign T799 = host_csr_req_fire & T800;
  assign T800 = host_csr_bits_rw ^ 1'h1;
  assign T801 = T804 & T802;
  assign T802 = T803 | host_csr_req_fire;
  assign T803 = reg_tohost == 64'h0;
  assign T804 = wen & T165;
  assign T805 = T810 | T973;
  assign T973 = {63'h0, T806};
  assign T806 = T167 ? reg_stats : 1'h0;
  assign T974 = reset ? 1'h0 : T807;
  assign T807 = T809 ? T808 : reg_stats;
  assign T808 = wdata[1'h0:1'h0];
  assign T809 = wen & T167;
  assign T810 = T812 | T975;
  assign T975 = {63'h0, T811};
  assign T811 = T169 ? io_host_id : 1'h0;
  assign T812 = T814 | T976;
  assign T976 = {63'h0, T813};
  assign T813 = T171 ? io_host_id : 1'h0;
  assign T814 = T816 | T815;
  assign T815 = T173 ? reg_mtimecmp : 64'h0;
  assign T816 = T818 | T817;
  assign T817 = T175 ? reg_mcause : 64'h0;
  assign T818 = T823 | T819;
  assign T819 = T177 ? T820 : 64'h0;
  assign T820 = {T821, reg_mbadaddr};
  assign T821 = 24'h0 - T977;
  assign T977 = {23'h0, T822};
  assign T822 = reg_mbadaddr[6'h27:6'h27];
  assign T823 = T828 | T824;
  assign T824 = T179 ? T825 : 64'h0;
  assign T825 = {T826, reg_mepc};
  assign T826 = 24'h0 - T978;
  assign T978 = {23'h0, T827};
  assign T827 = reg_mepc[6'h27:6'h27];
  assign T828 = T832 | T829;
  assign T829 = T181 ? reg_mscratch : 64'h0;
  assign T830 = T831 ? wdata : reg_mscratch;
  assign T831 = wen & T181;
  assign T832 = T842 | T979;
  assign T979 = {56'h0, T833};
  assign T833 = T183 ? T834 : 8'h0;
  assign T834 = T835;
  assign T835 = {T839, T836};
  assign T836 = {T838, T837};
  assign T837 = {reg_mie_ssip, reg_mie_usip};
  assign T980 = reset ? 1'h0 : reg_mie_usip;
  assign T838 = {reg_mie_msip, reg_mie_hsip};
  assign T981 = reset ? 1'h0 : reg_mie_hsip;
  assign T839 = {T841, T840};
  assign T840 = {reg_mie_stip, reg_mie_utip};
  assign T982 = reset ? 1'h0 : reg_mie_utip;
  assign T841 = {reg_mie_mtip, reg_mie_htip};
  assign T983 = reset ? 1'h0 : reg_mie_htip;
  assign T842 = T852 | T984;
  assign T984 = {56'h0, T843};
  assign T843 = T185 ? T844 : 8'h0;
  assign T844 = T845;
  assign T845 = {T849, T846};
  assign T846 = {T848, T847};
  assign T847 = {reg_mip_ssip, reg_mip_usip};
  assign T985 = reset ? 1'h0 : reg_mip_usip;
  assign T848 = {reg_mip_msip, reg_mip_hsip};
  assign T986 = reset ? 1'h0 : reg_mip_hsip;
  assign T849 = {T851, T850};
  assign T850 = {reg_mip_stip, reg_mip_utip};
  assign T987 = reset ? 1'h0 : reg_mip_utip;
  assign T851 = {reg_mip_mtip, reg_mip_htip};
  assign T988 = reset ? 1'h0 : reg_mip_htip;
  assign T852 = T854 | T989;
  assign T989 = {55'h0, T853};
  assign T853 = T187 ? 9'h100 : 9'h0;
  assign T854 = T855 | 64'h0;
  assign T855 = T856 | 64'h0;
  assign T856 = T858 | T857;
  assign T857 = T61 ? read_mstatus : 64'h0;
  assign T858 = T859 | T990;
  assign T990 = {63'h0, T194};
  assign T859 = T861 | T860;
  assign T860 = T196 ? 64'h8000000000041101 : 64'h0;
  assign T861 = T863 | T862;
  assign T862 = T198 ? read_time : 64'h0;
  assign T863 = T865 | T864;
  assign T864 = T200 ? read_time : 64'h0;
  assign T865 = T867 | T866;
  assign T866 = T202 ? read_time : 64'h0;
  assign T867 = T869 | T868;
  assign T868 = T204 ? read_time : 64'h0;
  assign T869 = T871 | T870;
  assign T870 = T206 ? read_time : 64'h0;
  assign T871 = T873 | T872;
  assign T872 = T208 ? T315 : 64'h0;
  assign T873 = 64'h0 | T874;
  assign T874 = T210 ? T315 : 64'h0;
  assign io_host_debug_stats_csr = reg_stats;
  assign io_host_ipi_rep_ready = 1'h1;
  assign io_host_ipi_req_bits = T991;
  assign T991 = io_rw_wdata[1'h0:1'h0];
  assign io_host_ipi_req_valid = T875;
  assign T875 = cpu_wen & T169;
  assign io_host_csr_resp_bits = host_csr_bits_data;
  assign io_host_csr_resp_valid = host_csr_rep_valid;
  assign T876 = T878 ? 1'h0 : T877;
  assign T877 = host_csr_req_fire ? 1'h1 : host_csr_rep_valid;
  assign T878 = io_host_csr_resp_ready & io_host_csr_resp_valid;
  assign io_host_csr_req_ready = T879;
  assign T879 = T881 & T880;
  assign T880 = host_csr_rep_valid ^ 1'h1;
  assign T881 = host_csr_req_valid ^ 1'h1;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "these conditions must be mutually exclusive");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      reg_mstatus_prv <= 2'h3;
    end else if(T90) begin
      reg_mstatus_prv <= T89;
    end else if(insn_redirect_trap) begin
      reg_mstatus_prv <= 2'h1;
    end else if(insn_ret) begin
      reg_mstatus_prv <= reg_mstatus_prv1;
    end else if(T27) begin
      reg_mstatus_prv <= 2'h3;
    end
    if(reset) begin
      reg_mstatus_prv1 <= 2'h3;
    end else if(T78) begin
      reg_mstatus_prv1 <= T883;
    end else if(T71) begin
      reg_mstatus_prv1 <= T70;
    end else if(insn_ret) begin
      reg_mstatus_prv1 <= reg_mstatus_prv2;
    end else if(T27) begin
      reg_mstatus_prv1 <= reg_mstatus_prv;
    end
    if(reset) begin
      reg_mstatus_prv2 <= 2'h0;
    end else if(T54) begin
      reg_mstatus_prv2 <= T37;
    end else if(insn_ret) begin
      reg_mstatus_prv2 <= 2'h0;
    end else if(T27) begin
      reg_mstatus_prv2 <= reg_mstatus_prv1;
    end
    if(host_csr_req_fire) begin
      host_csr_bits_data <= io_rw_rdata;
    end else if(T42) begin
      host_csr_bits_data <= io_host_csr_req_bits_data;
    end
    if(host_csr_req_fire) begin
      host_csr_req_valid <= 1'h0;
    end else if(T42) begin
      host_csr_req_valid <= 1'h1;
    end
    if(T42) begin
      host_csr_bits_addr <= io_host_csr_req_bits_addr;
    end
    if(T42) begin
      host_csr_bits_rw <= io_host_csr_req_bits_rw;
    end
    if(reset) begin
      reg_mstatus_ie <= 1'h0;
    end else if(T78) begin
      reg_mstatus_ie <= T243;
    end else if(T60) begin
      reg_mstatus_ie <= T242;
    end else if(insn_ret) begin
      reg_mstatus_ie <= reg_mstatus_ie1;
    end else if(T27) begin
      reg_mstatus_ie <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_ie1 <= 1'h0;
    end else if(T78) begin
      reg_mstatus_ie1 <= T241;
    end else if(T60) begin
      reg_mstatus_ie1 <= T240;
    end else if(insn_ret) begin
      reg_mstatus_ie1 <= reg_mstatus_ie2;
    end else if(T27) begin
      reg_mstatus_ie1 <= reg_mstatus_ie;
    end
    if(reset) begin
      reg_mstatus_ie2 <= 1'h0;
    end else if(T60) begin
      reg_mstatus_ie2 <= T239;
    end else if(insn_ret) begin
      reg_mstatus_ie2 <= 1'h1;
    end else if(T27) begin
      reg_mstatus_ie2 <= reg_mstatus_ie1;
    end
    if(reset) begin
      reg_mip_ssip <= 1'h0;
    end else if(T252) begin
      reg_mip_ssip <= T251;
    end else if(T250) begin
      reg_mip_ssip <= T249;
    end
    if(reset) begin
      reg_mie_ssip <= 1'h0;
    end else if(T258) begin
      reg_mie_ssip <= T257;
    end else if(T256) begin
      reg_mie_ssip <= T255;
    end
    if(reset) begin
      reg_mip_msip <= 1'h0;
    end else if(io_host_ipi_rep_valid) begin
      reg_mip_msip <= 1'h1;
    end else if(T250) begin
      reg_mip_msip <= T267;
    end
    if(reset) begin
      reg_mie_msip <= 1'h0;
    end else if(T256) begin
      reg_mie_msip <= T269;
    end
    if(reset) begin
      reg_mip_stip <= 1'h0;
    end else if(T250) begin
      reg_mip_stip <= T277;
    end
    if(reset) begin
      reg_mie_stip <= 1'h0;
    end else if(T258) begin
      reg_mie_stip <= T281;
    end else if(T256) begin
      reg_mie_stip <= T280;
    end
    if(reset) begin
      reg_mip_mtip <= 1'h0;
    end else if(T294) begin
      reg_mip_mtip <= 1'h0;
    end else if(T290) begin
      reg_mip_mtip <= 1'h1;
    end
    if(T292) begin
      read_time <= wdata;
    end
    if(T294) begin
      reg_mtimecmp <= wdata;
    end
    if(reset) begin
      reg_mie_mtip <= 1'h0;
    end else if(T256) begin
      reg_mie_mtip <= T296;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T304) begin
      reg_fromhost <= wdata;
    end
    reg_frm <= T896;
    if(reset) begin
      R316 <= 6'h0;
    end else begin
      R316 <= T317;
    end
    if(reset) begin
      R319 <= 58'h0;
    end else if(T322) begin
      R319 <= T321;
    end
    reg_sepc <= T902;
    reg_mepc <= T904;
    reg_stvec <= T906;
    if(T362) begin
      reg_sptbr <= T360;
    end
    if(reset) begin
      reg_mstatus_ie3 <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_prv3 <= 2'h0;
    end
    if(reset) begin
      reg_mstatus_fs <= 2'h0;
    end else if(T78) begin
      reg_mstatus_fs <= T371;
    end else if(T60) begin
      reg_mstatus_fs <= T370;
    end
    if(reset) begin
      reg_mstatus_xs <= 2'h0;
    end
    if(reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if(T78) begin
      reg_mstatus_mprv <= T380;
    end else if(T60) begin
      reg_mstatus_mprv <= T379;
    end else if(T27) begin
      reg_mstatus_mprv <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_vm <= 5'h0;
    end else if(T387) begin
      reg_mstatus_vm <= 5'h9;
    end else if(T384) begin
      reg_mstatus_vm <= 5'h0;
    end
    if(reset) begin
      reg_mstatus_zero1 <= 9'h0;
    end
    if(reset) begin
      reg_mstatus_sd_rv32 <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_zero2 <= 31'h0;
    end
    if(reset) begin
      reg_wfi <= 1'h0;
    end else if(some_interrupt_pending) begin
      reg_wfi <= 1'h0;
    end else if(insn_wfi) begin
      reg_wfi <= 1'h1;
    end
    if(insn_redirect_trap) begin
      reg_sbadaddr <= reg_mbadaddr;
    end
    if(T458) begin
      reg_mbadaddr <= T457;
    end else if(T449) begin
      reg_mbadaddr <= T441;
    end else if(T27) begin
      reg_mbadaddr <= io_pc;
    end
    if(insn_redirect_trap) begin
      reg_scause <= reg_mcause;
    end
    if(T474) begin
      reg_mcause <= T473;
    end else if(T472) begin
      reg_mcause <= T917;
    end else if(T470) begin
      reg_mcause <= 64'h3;
    end else if(T469) begin
      reg_mcause <= 64'h2;
    end else if(T27) begin
      reg_mcause <= io_cause;
    end
    if(T478) begin
      reg_sscratch <= wdata;
    end
    if(reset) begin
      R567 <= 6'h0;
    end else if(T571) begin
      R567 <= T569;
    end
    if(reset) begin
      R572 <= 58'h0;
    end else if(T575) begin
      R572 <= T574;
    end
    if(reset) begin
      R580 <= 6'h0;
    end else if(T584) begin
      R580 <= T582;
    end
    if(reset) begin
      R585 <= 58'h0;
    end else if(T588) begin
      R585 <= T587;
    end
    if(reset) begin
      R593 <= 6'h0;
    end else if(T597) begin
      R593 <= T595;
    end
    if(reset) begin
      R598 <= 58'h0;
    end else if(T601) begin
      R598 <= T600;
    end
    if(reset) begin
      R606 <= 6'h0;
    end else if(T610) begin
      R606 <= T608;
    end
    if(reset) begin
      R611 <= 58'h0;
    end else if(T614) begin
      R611 <= T613;
    end
    if(reset) begin
      R619 <= 6'h0;
    end else if(T623) begin
      R619 <= T621;
    end
    if(reset) begin
      R624 <= 58'h0;
    end else if(T627) begin
      R624 <= T626;
    end
    if(reset) begin
      R632 <= 6'h0;
    end else if(T636) begin
      R632 <= T634;
    end
    if(reset) begin
      R637 <= 58'h0;
    end else if(T640) begin
      R637 <= T639;
    end
    if(reset) begin
      R645 <= 6'h0;
    end else if(T649) begin
      R645 <= T647;
    end
    if(reset) begin
      R650 <= 58'h0;
    end else if(T653) begin
      R650 <= T652;
    end
    if(reset) begin
      R658 <= 6'h0;
    end else if(T662) begin
      R658 <= T660;
    end
    if(reset) begin
      R663 <= 58'h0;
    end else if(T666) begin
      R663 <= T665;
    end
    if(reset) begin
      R671 <= 6'h0;
    end else if(T675) begin
      R671 <= T673;
    end
    if(reset) begin
      R676 <= 58'h0;
    end else if(T679) begin
      R676 <= T678;
    end
    if(reset) begin
      R684 <= 6'h0;
    end else if(T688) begin
      R684 <= T686;
    end
    if(reset) begin
      R689 <= 58'h0;
    end else if(T692) begin
      R689 <= T691;
    end
    if(reset) begin
      R697 <= 6'h0;
    end else if(T701) begin
      R697 <= T699;
    end
    if(reset) begin
      R702 <= 58'h0;
    end else if(T705) begin
      R702 <= T704;
    end
    if(reset) begin
      R710 <= 6'h0;
    end else if(T714) begin
      R710 <= T712;
    end
    if(reset) begin
      R715 <= 58'h0;
    end else if(T718) begin
      R715 <= T717;
    end
    if(reset) begin
      R723 <= 6'h0;
    end else if(T727) begin
      R723 <= T725;
    end
    if(reset) begin
      R728 <= 58'h0;
    end else if(T731) begin
      R728 <= T730;
    end
    if(reset) begin
      R736 <= 6'h0;
    end else if(T740) begin
      R736 <= T738;
    end
    if(reset) begin
      R741 <= 58'h0;
    end else if(T744) begin
      R741 <= T743;
    end
    if(reset) begin
      R749 <= 6'h0;
    end else if(T753) begin
      R749 <= T751;
    end
    if(reset) begin
      R754 <= 58'h0;
    end else if(T757) begin
      R754 <= T756;
    end
    if(reset) begin
      R762 <= 6'h0;
    end else if(T766) begin
      R762 <= T764;
    end
    if(reset) begin
      R767 <= 58'h0;
    end else if(T770) begin
      R767 <= T769;
    end
    if(reset) begin
      R775 <= 6'h0;
    end else if(T782) begin
      R775 <= T781;
    end else if(T780) begin
      R775 <= T778;
    end
    if(reset) begin
      R783 <= 58'h0;
    end else if(T782) begin
      R783 <= T789;
    end else if(T787) begin
      R783 <= T786;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T801) begin
      reg_tohost <= wdata;
    end else if(T798) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T809) begin
      reg_stats <= T808;
    end
    if(T831) begin
      reg_mscratch <= wdata;
    end
    if(reset) begin
      reg_mie_usip <= 1'h0;
    end
    if(reset) begin
      reg_mie_hsip <= 1'h0;
    end
    if(reset) begin
      reg_mie_utip <= 1'h0;
    end
    if(reset) begin
      reg_mie_htip <= 1'h0;
    end
    if(reset) begin
      reg_mip_usip <= 1'h0;
    end
    if(reset) begin
      reg_mip_hsip <= 1'h0;
    end
    if(reset) begin
      reg_mip_utip <= 1'h0;
    end
    if(reset) begin
      reg_mip_htip <= 1'h0;
    end
    if(T878) begin
      host_csr_rep_valid <= 1'h0;
    end else if(host_csr_req_fire) begin
      host_csr_rep_valid <= 1'h1;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out
);

  wire[63:0] sum;
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[31:0] T5;
  wire[63:0] out64;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T136;
  wire cmp;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[63:0] T25;
  wire T26;
  wire[63:0] T27;
  wire T28;
  wire[63:0] T29;
  wire T30;
  wire[63:0] shout_l;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[62:0] T33;
  wire[63:0] T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire[61:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[59:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  wire[63:0] T44;
  wire[55:0] T45;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[47:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[31:0] T53;
  wire[63:0] T54;
  wire[63:0] T137;
  wire[31:0] T55;
  wire[63:0] T56;
  wire[63:0] T138;
  wire[47:0] T57;
  wire[63:0] T58;
  wire[63:0] T139;
  wire[55:0] T59;
  wire[63:0] T60;
  wire[63:0] T140;
  wire[59:0] T61;
  wire[63:0] T62;
  wire[63:0] T141;
  wire[61:0] T63;
  wire[63:0] T64;
  wire[63:0] T142;
  wire[62:0] T65;
  wire T66;
  wire[63:0] shout_r;
  wire[64:0] T67;
  wire[5:0] shamt;
  wire[5:0] T68;
  wire[4:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[64:0] T74;
  wire[64:0] T75;
  wire[63:0] shin;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[63:0] T78;
  wire[62:0] T79;
  wire[63:0] T80;
  wire[63:0] T81;
  wire[63:0] T82;
  wire[61:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[59:0] T87;
  wire[63:0] T88;
  wire[63:0] T89;
  wire[63:0] T90;
  wire[55:0] T91;
  wire[63:0] T92;
  wire[63:0] T93;
  wire[63:0] T94;
  wire[47:0] T95;
  wire[63:0] T96;
  wire[63:0] T97;
  wire[63:0] T98;
  wire[31:0] T99;
  wire[63:0] T100;
  wire[63:0] T143;
  wire[31:0] T101;
  wire[63:0] T102;
  wire[63:0] T144;
  wire[47:0] T103;
  wire[63:0] T104;
  wire[63:0] T145;
  wire[55:0] T105;
  wire[63:0] T106;
  wire[63:0] T146;
  wire[59:0] T107;
  wire[63:0] T108;
  wire[63:0] T147;
  wire[61:0] T109;
  wire[63:0] T110;
  wire[63:0] T148;
  wire[62:0] T111;
  wire[63:0] shin_r;
  wire[31:0] T112;
  wire[31:0] shin_hi;
  wire[31:0] shin_hi_32;
  wire[31:0] T113;
  wire[31:0] T149;
  wire T114;
  wire T115;
  wire[31:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire[31:0] out_hi;
  wire[31:0] T131;
  wire[31:0] T150;
  wire T132;
  wire[31:0] T133;
  wire T134;
  wire T135;


  assign io_adder_out = sum;
  assign sum = io_in1 + T0;
  assign T0 = T2 ? T1 : io_in2;
  assign T1 = 64'h0 - io_in2;
  assign T2 = io_fn[2'h3:2'h3];
  assign io_out = T3;
  assign T3 = T4;
  assign T4 = {out_hi, T5};
  assign T5 = out64[5'h1f:1'h0];
  assign out64 = T128 ? sum : T6;
  assign T6 = T125 ? shout_r : T7;
  assign T7 = T66 ? shout_l : T8;
  assign T8 = T30 ? T29 : T9;
  assign T9 = T28 ? T27 : T10;
  assign T10 = T26 ? T25 : T136;
  assign T136 = {63'h0, cmp};
  assign cmp = T24 ^ T11;
  assign T11 = T22 ? T21 : T12;
  assign T12 = T18 ? T17 : T13;
  assign T13 = T16 ? T15 : T14;
  assign T14 = io_in1[6'h3f:6'h3f];
  assign T15 = io_in2[6'h3f:6'h3f];
  assign T16 = io_fn[1'h1:1'h1];
  assign T17 = sum[6'h3f:6'h3f];
  assign T18 = T20 == T19;
  assign T19 = io_in2[6'h3f:6'h3f];
  assign T20 = io_in1[6'h3f:6'h3f];
  assign T21 = sum == 64'h0;
  assign T22 = T23 ^ 1'h1;
  assign T23 = io_fn[2'h2:2'h2];
  assign T24 = io_fn[1'h0:1'h0];
  assign T25 = io_in1 ^ io_in2;
  assign T26 = io_fn == 4'h4;
  assign T27 = io_in1 | io_in2;
  assign T28 = io_fn == 4'h6;
  assign T29 = io_in1 & io_in2;
  assign T30 = io_fn == 4'h7;
  assign shout_l = T64 | T31;
  assign T31 = T32 & 64'haaaaaaaaaaaaaaaa;
  assign T32 = T33 << 1'h1;
  assign T33 = T34[6'h3e:1'h0];
  assign T34 = T62 | T35;
  assign T35 = T36 & 64'hcccccccccccccccc;
  assign T36 = T37 << 2'h2;
  assign T37 = T38[6'h3d:1'h0];
  assign T38 = T60 | T39;
  assign T39 = T40 & 64'hf0f0f0f0f0f0f0f0;
  assign T40 = T41 << 3'h4;
  assign T41 = T42[6'h3b:1'h0];
  assign T42 = T58 | T43;
  assign T43 = T44 & 64'hff00ff00ff00ff00;
  assign T44 = T45 << 4'h8;
  assign T45 = T46[6'h37:1'h0];
  assign T46 = T56 | T47;
  assign T47 = T48 & 64'hffff0000ffff0000;
  assign T48 = T49 << 5'h10;
  assign T49 = T50[6'h2f:1'h0];
  assign T50 = T54 | T51;
  assign T51 = T52 & 64'hffffffff00000000;
  assign T52 = T53 << 6'h20;
  assign T53 = shout_r[5'h1f:1'h0];
  assign T54 = T137 & 64'hffffffff;
  assign T137 = {32'h0, T55};
  assign T55 = shout_r >> 6'h20;
  assign T56 = T138 & 64'hffff0000ffff;
  assign T138 = {16'h0, T57};
  assign T57 = T50 >> 5'h10;
  assign T58 = T139 & 64'hff00ff00ff00ff;
  assign T139 = {8'h0, T59};
  assign T59 = T46 >> 4'h8;
  assign T60 = T140 & 64'hf0f0f0f0f0f0f0f;
  assign T140 = {4'h0, T61};
  assign T61 = T42 >> 3'h4;
  assign T62 = T141 & 64'h3333333333333333;
  assign T141 = {2'h0, T63};
  assign T63 = T38 >> 2'h2;
  assign T64 = T142 & 64'h5555555555555555;
  assign T142 = {1'h0, T65};
  assign T65 = T34 >> 1'h1;
  assign T66 = io_fn == 4'h1;
  assign shout_r = T67[6'h3f:1'h0];
  assign T67 = $signed(T74) >>> shamt;
  assign shamt = T68;
  assign T68 = {T70, T69};
  assign T69 = io_in2[3'h4:1'h0];
  assign T70 = T73 & T71;
  assign T71 = 1'h1 == T72;
  assign T72 = io_dw & 1'h1;
  assign T73 = io_in2[3'h5:3'h5];
  assign T74 = T75;
  assign T75 = {T122, shin};
  assign shin = T119 ? shin_r : T76;
  assign T76 = T110 | T77;
  assign T77 = T78 & 64'haaaaaaaaaaaaaaaa;
  assign T78 = T79 << 1'h1;
  assign T79 = T80[6'h3e:1'h0];
  assign T80 = T108 | T81;
  assign T81 = T82 & 64'hcccccccccccccccc;
  assign T82 = T83 << 2'h2;
  assign T83 = T84[6'h3d:1'h0];
  assign T84 = T106 | T85;
  assign T85 = T86 & 64'hf0f0f0f0f0f0f0f0;
  assign T86 = T87 << 3'h4;
  assign T87 = T88[6'h3b:1'h0];
  assign T88 = T104 | T89;
  assign T89 = T90 & 64'hff00ff00ff00ff00;
  assign T90 = T91 << 4'h8;
  assign T91 = T92[6'h37:1'h0];
  assign T92 = T102 | T93;
  assign T93 = T94 & 64'hffff0000ffff0000;
  assign T94 = T95 << 5'h10;
  assign T95 = T96[6'h2f:1'h0];
  assign T96 = T100 | T97;
  assign T97 = T98 & 64'hffffffff00000000;
  assign T98 = T99 << 6'h20;
  assign T99 = shin_r[5'h1f:1'h0];
  assign T100 = T143 & 64'hffffffff;
  assign T143 = {32'h0, T101};
  assign T101 = shin_r >> 6'h20;
  assign T102 = T144 & 64'hffff0000ffff;
  assign T144 = {16'h0, T103};
  assign T103 = T96 >> 5'h10;
  assign T104 = T145 & 64'hff00ff00ff00ff;
  assign T145 = {8'h0, T105};
  assign T105 = T92 >> 4'h8;
  assign T106 = T146 & 64'hf0f0f0f0f0f0f0f;
  assign T146 = {4'h0, T107};
  assign T107 = T88 >> 3'h4;
  assign T108 = T147 & 64'h3333333333333333;
  assign T147 = {2'h0, T109};
  assign T109 = T84 >> 2'h2;
  assign T110 = T148 & 64'h5555555555555555;
  assign T148 = {1'h0, T111};
  assign T111 = T80 >> 1'h1;
  assign shin_r = {shin_hi, T112};
  assign T112 = io_in1[5'h1f:1'h0];
  assign shin_hi = T117 ? T116 : shin_hi_32;
  assign shin_hi_32 = T115 ? T113 : 32'h0;
  assign T113 = 32'h0 - T149;
  assign T149 = {31'h0, T114};
  assign T114 = io_in1[5'h1f:5'h1f];
  assign T115 = io_fn[2'h3:2'h3];
  assign T116 = io_in1[6'h3f:6'h20];
  assign T117 = 1'h1 == T118;
  assign T118 = io_dw & 1'h1;
  assign T119 = T121 | T120;
  assign T120 = io_fn == 4'hb;
  assign T121 = io_fn == 4'h5;
  assign T122 = T124 & T123;
  assign T123 = shin[6'h3f:6'h3f];
  assign T124 = io_fn[2'h3:2'h3];
  assign T125 = T127 | T126;
  assign T126 = io_fn == 4'hb;
  assign T127 = io_fn == 4'h5;
  assign T128 = T130 | T129;
  assign T129 = io_fn == 4'ha;
  assign T130 = io_fn == 4'h0;
  assign out_hi = T134 ? T133 : T131;
  assign T131 = 32'h0 - T150;
  assign T150 = {31'h0, T132};
  assign T132 = out64[5'h1f:5'h1f];
  assign T133 = out64[6'h3f:6'h20];
  assign T134 = 1'h1 == T135;
  assign T135 = io_dw & 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T10;
  wire[129:0] T188;
  wire[63:0] negated_remainder;
  wire[63:0] T126;
  wire T11;
  wire T12;
  reg  isMul;
  wire T13;
  wire cmdMul;
  wire T14;
  wire T15;
  wire[3:0] T16;
  wire T17;
  wire[3:0] T18;
  wire T19;
  wire T20;
  reg [2:0] state;
  wire[2:0] T189;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  reg  neg_out;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  isHi;
  wire T34;
  wire cmdHi;
  wire T35;
  wire T36;
  wire T37;
  wire[3:0] T38;
  wire T39;
  wire[3:0] T40;
  wire T41;
  wire T42;
  wire less;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T43;
  wire[64:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[64:0] T48;
  wire[63:0] rhs_in;
  wire[31:0] T49;
  wire[31:0] T50;
  wire[31:0] T51;
  wire[31:0] T190;
  wire[31:0] T52;
  wire T53;
  wire T54;
  wire rhs_sign;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire rhsSigned;
  wire T60;
  wire T61;
  wire[3:0] T62;
  wire[64:0] T63;
  wire T64;
  reg [6:0] count;
  wire[6:0] T65;
  wire[6:0] T66;
  wire[6:0] T67;
  wire[6:0] T68;
  wire[6:0] T69;
  wire[6:0] T70;
  wire[6:0] T191;
  wire[5:0] T71;
  wire[5:0] T72;
  wire[5:0] T73;
  wire[5:0] T192;
  wire[5:0] T193;
  wire[5:0] T194;
  wire[5:0] T195;
  wire[5:0] T196;
  wire[5:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[5:0] T200;
  wire[5:0] T201;
  wire[5:0] T202;
  wire[5:0] T203;
  wire[5:0] T204;
  wire[5:0] T205;
  wire[5:0] T206;
  wire[5:0] T207;
  wire[5:0] T208;
  wire[5:0] T209;
  wire[5:0] T210;
  wire[5:0] T211;
  wire[5:0] T212;
  wire[5:0] T213;
  wire[5:0] T214;
  wire[5:0] T215;
  wire[5:0] T216;
  wire[5:0] T217;
  wire[5:0] T218;
  wire[5:0] T219;
  wire[5:0] T220;
  wire[5:0] T221;
  wire[5:0] T222;
  wire[5:0] T223;
  wire[4:0] T224;
  wire[4:0] T225;
  wire[4:0] T226;
  wire[4:0] T227;
  wire[4:0] T228;
  wire[4:0] T229;
  wire[4:0] T230;
  wire[4:0] T231;
  wire[4:0] T232;
  wire[4:0] T233;
  wire[4:0] T234;
  wire[4:0] T235;
  wire[4:0] T236;
  wire[4:0] T237;
  wire[4:0] T238;
  wire[4:0] T239;
  wire[3:0] T240;
  wire[3:0] T241;
  wire[3:0] T242;
  wire[3:0] T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[3:0] T246;
  wire[3:0] T247;
  wire[2:0] T248;
  wire[2:0] T249;
  wire[2:0] T250;
  wire[2:0] T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire T254;
  wire[63:0] T75;
  wire[63:0] T76;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire[5:0] T77;
  wire[5:0] T317;
  wire[5:0] T318;
  wire[5:0] T319;
  wire[5:0] T320;
  wire[5:0] T321;
  wire[5:0] T322;
  wire[5:0] T323;
  wire[5:0] T324;
  wire[5:0] T325;
  wire[5:0] T326;
  wire[5:0] T327;
  wire[5:0] T328;
  wire[5:0] T329;
  wire[5:0] T330;
  wire[5:0] T331;
  wire[5:0] T332;
  wire[5:0] T333;
  wire[5:0] T334;
  wire[5:0] T335;
  wire[5:0] T336;
  wire[5:0] T337;
  wire[5:0] T338;
  wire[5:0] T339;
  wire[5:0] T340;
  wire[5:0] T341;
  wire[5:0] T342;
  wire[5:0] T343;
  wire[5:0] T344;
  wire[5:0] T345;
  wire[5:0] T346;
  wire[5:0] T347;
  wire[5:0] T348;
  wire[4:0] T349;
  wire[4:0] T350;
  wire[4:0] T351;
  wire[4:0] T352;
  wire[4:0] T353;
  wire[4:0] T354;
  wire[4:0] T355;
  wire[4:0] T356;
  wire[4:0] T357;
  wire[4:0] T358;
  wire[4:0] T359;
  wire[4:0] T360;
  wire[4:0] T361;
  wire[4:0] T362;
  wire[4:0] T363;
  wire[4:0] T364;
  wire[3:0] T365;
  wire[3:0] T366;
  wire[3:0] T367;
  wire[3:0] T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire[3:0] T371;
  wire[3:0] T372;
  wire[2:0] T373;
  wire[2:0] T374;
  wire[2:0] T375;
  wire[2:0] T376;
  wire[1:0] T377;
  wire[1:0] T378;
  wire T379;
  wire[63:0] T79;
  wire[63:0] T80;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire lhs_sign;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire lhsSigned;
  wire T90;
  wire T91;
  wire[3:0] T92;
  wire T93;
  wire T94;
  wire[2:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire[63:0] T101;
  wire[63:0] T102;
  wire[63:0] T103;
  wire[64:0] T104;
  wire[5:0] T105;
  wire[10:0] T106;
  wire[63:0] T107;
  wire[128:0] T108;
  wire[63:0] T109;
  wire[64:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[2:0] T116;
  wire[2:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire T123;
  wire T124;
  wire T125;
  wire[129:0] T442;
  wire T127;
  wire[129:0] T443;
  wire[63:0] T128;
  wire T129;
  wire[129:0] T130;
  wire[64:0] T131;
  wire[63:0] T132;
  wire[128:0] T133;
  wire[63:0] T134;
  wire[128:0] T135;
  wire[128:0] T136;
  wire[128:0] T137;
  wire[55:0] T138;
  wire[72:0] T139;
  wire[72:0] T444;
  wire[64:0] T140;
  wire[64:0] T141;
  wire[7:0] T445;
  wire T446;
  wire[72:0] T142;
  wire[8:0] T143;
  wire[8:0] T144;
  wire[7:0] T145;
  wire[64:0] T146;
  wire[128:0] T147;
  wire[5:0] T148;
  wire[10:0] T149;
  wire[10:0] T150;
  wire[64:0] T151;
  wire[64:0] T152;
  wire T153;
  wire T154;
  wire[129:0] T447;
  wire[128:0] T155;
  wire[64:0] T156;
  wire T157;
  wire[63:0] T158;
  wire[63:0] T159;
  wire[63:0] T160;
  wire[63:0] T161;
  wire T162;
  wire T163;
  wire T164;
  wire[129:0] T448;
  wire[126:0] T165;
  wire[63:0] T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[129:0] T449;
  wire[63:0] lhs_in;
  wire[31:0] T173;
  wire[31:0] T174;
  wire[31:0] T175;
  wire[31:0] T450;
  wire[31:0] T176;
  wire T177;
  wire T178;
  wire[63:0] T179;
  wire[31:0] T180;
  wire[31:0] T181;
  wire[31:0] T451;
  wire T182;
  wire T183;
  wire T184;
  reg  req_dw;
  wire T185;
  wire T186;
  wire T187;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T183 ? T179 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T449 : T5;
  assign T5 = T167 ? T448 : T6;
  assign T6 = T162 ? T447 : T7;
  assign T7 = T153 ? T130 : T8;
  assign T8 = T129 ? T443 : T9;
  assign T9 = T127 ? T442 : T10;
  assign T10 = T11 ? T188 : remainder;
  assign T188 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T126;
  assign T126 = remainder[6'h3f:1'h0];
  assign T11 = T20 & T12;
  assign T12 = T19 | isMul;
  assign T13 = T1 ? cmdMul : isMul;
  assign cmdMul = T14;
  assign T14 = T17 | T15;
  assign T15 = T16 == 4'h8;
  assign T16 = io_req_bits_fn & 4'h8;
  assign T17 = T18 == 4'h0;
  assign T18 = io_req_bits_fn & 4'h4;
  assign T19 = remainder[6'h3f:6'h3f];
  assign T20 = state == 3'h1;
  assign T189 = reset ? 3'h0 : T21;
  assign T21 = T1 ? T122 : T22;
  assign T22 = T120 ? 3'h0 : T23;
  assign T23 = T118 ? T116 : T24;
  assign T24 = T96 ? T95 : T25;
  assign T25 = T129 ? T28 : T26;
  assign T26 = T127 ? 3'h5 : T27;
  assign T27 = T20 ? 3'h2 : state;
  assign T28 = neg_out ? 3'h4 : 3'h5;
  assign T29 = T1 ? T82 : T30;
  assign T30 = T31 ? 1'h0 : neg_out;
  assign T31 = T162 & T32;
  assign T32 = T41 & T33;
  assign T33 = isHi ^ 1'h1;
  assign T34 = T1 ? cmdHi : isHi;
  assign cmdHi = T35;
  assign T35 = T36 | T15;
  assign T36 = T39 | T37;
  assign T37 = T38 == 4'h2;
  assign T38 = io_req_bits_fn & 4'h2;
  assign T39 = T40 == 4'h1;
  assign T40 = io_req_bits_fn & 4'h5;
  assign T41 = T64 & T42;
  assign T42 = less ^ 1'h1;
  assign less = subtractor[7'h40:7'h40];
  assign subtractor = T63 - divisor;
  assign T43 = T1 ? T48 : T44;
  assign T44 = T45 ? subtractor : divisor;
  assign T45 = T20 & T46;
  assign T46 = T47 | isMul;
  assign T47 = divisor[6'h3f:6'h3f];
  assign T48 = {rhs_sign, rhs_in};
  assign rhs_in = {T50, T49};
  assign T49 = io_req_bits_in2[5'h1f:1'h0];
  assign T50 = T53 ? T52 : T51;
  assign T51 = 32'h0 - T190;
  assign T190 = {31'h0, rhs_sign};
  assign T52 = io_req_bits_in2[6'h3f:6'h20];
  assign T53 = 1'h1 == T54;
  assign T54 = io_req_bits_dw & 1'h1;
  assign rhs_sign = rhsSigned & T55;
  assign T55 = T58 ? T57 : T56;
  assign T56 = io_req_bits_in2[5'h1f:5'h1f];
  assign T57 = io_req_bits_in2[6'h3f:6'h3f];
  assign T58 = 1'h1 == T59;
  assign T59 = io_req_bits_dw & 1'h1;
  assign rhsSigned = T60;
  assign T60 = T61 | T17;
  assign T61 = T62 == 4'h0;
  assign T62 = io_req_bits_fn & 4'h9;
  assign T63 = remainder[8'h80:7'h40];
  assign T64 = count == 7'h0;
  assign T65 = T1 ? 7'h0 : T66;
  assign T66 = T167 ? T191 : T67;
  assign T67 = T162 ? T70 : T68;
  assign T68 = T153 ? T69 : count;
  assign T69 = count + 7'h1;
  assign T70 = count + 7'h1;
  assign T191 = {1'h0, T71};
  assign T71 = T81 ? 6'h3f : T72;
  assign T72 = T73[3'h5:1'h0];
  assign T73 = T77 - T192;
  assign T192 = T316 ? 6'h3f : T193;
  assign T193 = T315 ? 6'h3e : T194;
  assign T194 = T314 ? 6'h3d : T195;
  assign T195 = T313 ? 6'h3c : T196;
  assign T196 = T312 ? 6'h3b : T197;
  assign T197 = T311 ? 6'h3a : T198;
  assign T198 = T310 ? 6'h39 : T199;
  assign T199 = T309 ? 6'h38 : T200;
  assign T200 = T308 ? 6'h37 : T201;
  assign T201 = T307 ? 6'h36 : T202;
  assign T202 = T306 ? 6'h35 : T203;
  assign T203 = T305 ? 6'h34 : T204;
  assign T204 = T304 ? 6'h33 : T205;
  assign T205 = T303 ? 6'h32 : T206;
  assign T206 = T302 ? 6'h31 : T207;
  assign T207 = T301 ? 6'h30 : T208;
  assign T208 = T300 ? 6'h2f : T209;
  assign T209 = T299 ? 6'h2e : T210;
  assign T210 = T298 ? 6'h2d : T211;
  assign T211 = T297 ? 6'h2c : T212;
  assign T212 = T296 ? 6'h2b : T213;
  assign T213 = T295 ? 6'h2a : T214;
  assign T214 = T294 ? 6'h29 : T215;
  assign T215 = T293 ? 6'h28 : T216;
  assign T216 = T292 ? 6'h27 : T217;
  assign T217 = T291 ? 6'h26 : T218;
  assign T218 = T290 ? 6'h25 : T219;
  assign T219 = T289 ? 6'h24 : T220;
  assign T220 = T288 ? 6'h23 : T221;
  assign T221 = T287 ? 6'h22 : T222;
  assign T222 = T286 ? 6'h21 : T223;
  assign T223 = T285 ? 6'h20 : T224;
  assign T224 = T284 ? 5'h1f : T225;
  assign T225 = T283 ? 5'h1e : T226;
  assign T226 = T282 ? 5'h1d : T227;
  assign T227 = T281 ? 5'h1c : T228;
  assign T228 = T280 ? 5'h1b : T229;
  assign T229 = T279 ? 5'h1a : T230;
  assign T230 = T278 ? 5'h19 : T231;
  assign T231 = T277 ? 5'h18 : T232;
  assign T232 = T276 ? 5'h17 : T233;
  assign T233 = T275 ? 5'h16 : T234;
  assign T234 = T274 ? 5'h15 : T235;
  assign T235 = T273 ? 5'h14 : T236;
  assign T236 = T272 ? 5'h13 : T237;
  assign T237 = T271 ? 5'h12 : T238;
  assign T238 = T270 ? 5'h11 : T239;
  assign T239 = T269 ? 5'h10 : T240;
  assign T240 = T268 ? 4'hf : T241;
  assign T241 = T267 ? 4'he : T242;
  assign T242 = T266 ? 4'hd : T243;
  assign T243 = T265 ? 4'hc : T244;
  assign T244 = T264 ? 4'hb : T245;
  assign T245 = T263 ? 4'ha : T246;
  assign T246 = T262 ? 4'h9 : T247;
  assign T247 = T261 ? 4'h8 : T248;
  assign T248 = T260 ? 3'h7 : T249;
  assign T249 = T259 ? 3'h6 : T250;
  assign T250 = T258 ? 3'h5 : T251;
  assign T251 = T257 ? 3'h4 : T252;
  assign T252 = T256 ? 2'h3 : T253;
  assign T253 = T255 ? 2'h2 : T254;
  assign T254 = T75[1'h1:1'h1];
  assign T75 = T76[6'h3f:1'h0];
  assign T76 = remainder[6'h3f:1'h0];
  assign T255 = T75[2'h2:2'h2];
  assign T256 = T75[2'h3:2'h3];
  assign T257 = T75[3'h4:3'h4];
  assign T258 = T75[3'h5:3'h5];
  assign T259 = T75[3'h6:3'h6];
  assign T260 = T75[3'h7:3'h7];
  assign T261 = T75[4'h8:4'h8];
  assign T262 = T75[4'h9:4'h9];
  assign T263 = T75[4'ha:4'ha];
  assign T264 = T75[4'hb:4'hb];
  assign T265 = T75[4'hc:4'hc];
  assign T266 = T75[4'hd:4'hd];
  assign T267 = T75[4'he:4'he];
  assign T268 = T75[4'hf:4'hf];
  assign T269 = T75[5'h10:5'h10];
  assign T270 = T75[5'h11:5'h11];
  assign T271 = T75[5'h12:5'h12];
  assign T272 = T75[5'h13:5'h13];
  assign T273 = T75[5'h14:5'h14];
  assign T274 = T75[5'h15:5'h15];
  assign T275 = T75[5'h16:5'h16];
  assign T276 = T75[5'h17:5'h17];
  assign T277 = T75[5'h18:5'h18];
  assign T278 = T75[5'h19:5'h19];
  assign T279 = T75[5'h1a:5'h1a];
  assign T280 = T75[5'h1b:5'h1b];
  assign T281 = T75[5'h1c:5'h1c];
  assign T282 = T75[5'h1d:5'h1d];
  assign T283 = T75[5'h1e:5'h1e];
  assign T284 = T75[5'h1f:5'h1f];
  assign T285 = T75[6'h20:6'h20];
  assign T286 = T75[6'h21:6'h21];
  assign T287 = T75[6'h22:6'h22];
  assign T288 = T75[6'h23:6'h23];
  assign T289 = T75[6'h24:6'h24];
  assign T290 = T75[6'h25:6'h25];
  assign T291 = T75[6'h26:6'h26];
  assign T292 = T75[6'h27:6'h27];
  assign T293 = T75[6'h28:6'h28];
  assign T294 = T75[6'h29:6'h29];
  assign T295 = T75[6'h2a:6'h2a];
  assign T296 = T75[6'h2b:6'h2b];
  assign T297 = T75[6'h2c:6'h2c];
  assign T298 = T75[6'h2d:6'h2d];
  assign T299 = T75[6'h2e:6'h2e];
  assign T300 = T75[6'h2f:6'h2f];
  assign T301 = T75[6'h30:6'h30];
  assign T302 = T75[6'h31:6'h31];
  assign T303 = T75[6'h32:6'h32];
  assign T304 = T75[6'h33:6'h33];
  assign T305 = T75[6'h34:6'h34];
  assign T306 = T75[6'h35:6'h35];
  assign T307 = T75[6'h36:6'h36];
  assign T308 = T75[6'h37:6'h37];
  assign T309 = T75[6'h38:6'h38];
  assign T310 = T75[6'h39:6'h39];
  assign T311 = T75[6'h3a:6'h3a];
  assign T312 = T75[6'h3b:6'h3b];
  assign T313 = T75[6'h3c:6'h3c];
  assign T314 = T75[6'h3d:6'h3d];
  assign T315 = T75[6'h3e:6'h3e];
  assign T316 = T75[6'h3f:6'h3f];
  assign T77 = 6'h3f + T317;
  assign T317 = T441 ? 6'h3f : T318;
  assign T318 = T440 ? 6'h3e : T319;
  assign T319 = T439 ? 6'h3d : T320;
  assign T320 = T438 ? 6'h3c : T321;
  assign T321 = T437 ? 6'h3b : T322;
  assign T322 = T436 ? 6'h3a : T323;
  assign T323 = T435 ? 6'h39 : T324;
  assign T324 = T434 ? 6'h38 : T325;
  assign T325 = T433 ? 6'h37 : T326;
  assign T326 = T432 ? 6'h36 : T327;
  assign T327 = T431 ? 6'h35 : T328;
  assign T328 = T430 ? 6'h34 : T329;
  assign T329 = T429 ? 6'h33 : T330;
  assign T330 = T428 ? 6'h32 : T331;
  assign T331 = T427 ? 6'h31 : T332;
  assign T332 = T426 ? 6'h30 : T333;
  assign T333 = T425 ? 6'h2f : T334;
  assign T334 = T424 ? 6'h2e : T335;
  assign T335 = T423 ? 6'h2d : T336;
  assign T336 = T422 ? 6'h2c : T337;
  assign T337 = T421 ? 6'h2b : T338;
  assign T338 = T420 ? 6'h2a : T339;
  assign T339 = T419 ? 6'h29 : T340;
  assign T340 = T418 ? 6'h28 : T341;
  assign T341 = T417 ? 6'h27 : T342;
  assign T342 = T416 ? 6'h26 : T343;
  assign T343 = T415 ? 6'h25 : T344;
  assign T344 = T414 ? 6'h24 : T345;
  assign T345 = T413 ? 6'h23 : T346;
  assign T346 = T412 ? 6'h22 : T347;
  assign T347 = T411 ? 6'h21 : T348;
  assign T348 = T410 ? 6'h20 : T349;
  assign T349 = T409 ? 5'h1f : T350;
  assign T350 = T408 ? 5'h1e : T351;
  assign T351 = T407 ? 5'h1d : T352;
  assign T352 = T406 ? 5'h1c : T353;
  assign T353 = T405 ? 5'h1b : T354;
  assign T354 = T404 ? 5'h1a : T355;
  assign T355 = T403 ? 5'h19 : T356;
  assign T356 = T402 ? 5'h18 : T357;
  assign T357 = T401 ? 5'h17 : T358;
  assign T358 = T400 ? 5'h16 : T359;
  assign T359 = T399 ? 5'h15 : T360;
  assign T360 = T398 ? 5'h14 : T361;
  assign T361 = T397 ? 5'h13 : T362;
  assign T362 = T396 ? 5'h12 : T363;
  assign T363 = T395 ? 5'h11 : T364;
  assign T364 = T394 ? 5'h10 : T365;
  assign T365 = T393 ? 4'hf : T366;
  assign T366 = T392 ? 4'he : T367;
  assign T367 = T391 ? 4'hd : T368;
  assign T368 = T390 ? 4'hc : T369;
  assign T369 = T389 ? 4'hb : T370;
  assign T370 = T388 ? 4'ha : T371;
  assign T371 = T387 ? 4'h9 : T372;
  assign T372 = T386 ? 4'h8 : T373;
  assign T373 = T385 ? 3'h7 : T374;
  assign T374 = T384 ? 3'h6 : T375;
  assign T375 = T383 ? 3'h5 : T376;
  assign T376 = T382 ? 3'h4 : T377;
  assign T377 = T381 ? 2'h3 : T378;
  assign T378 = T380 ? 2'h2 : T379;
  assign T379 = T79[1'h1:1'h1];
  assign T79 = T80[6'h3f:1'h0];
  assign T80 = divisor[6'h3f:1'h0];
  assign T380 = T79[2'h2:2'h2];
  assign T381 = T79[2'h3:2'h3];
  assign T382 = T79[3'h4:3'h4];
  assign T383 = T79[3'h5:3'h5];
  assign T384 = T79[3'h6:3'h6];
  assign T385 = T79[3'h7:3'h7];
  assign T386 = T79[4'h8:4'h8];
  assign T387 = T79[4'h9:4'h9];
  assign T388 = T79[4'ha:4'ha];
  assign T389 = T79[4'hb:4'hb];
  assign T390 = T79[4'hc:4'hc];
  assign T391 = T79[4'hd:4'hd];
  assign T392 = T79[4'he:4'he];
  assign T393 = T79[4'hf:4'hf];
  assign T394 = T79[5'h10:5'h10];
  assign T395 = T79[5'h11:5'h11];
  assign T396 = T79[5'h12:5'h12];
  assign T397 = T79[5'h13:5'h13];
  assign T398 = T79[5'h14:5'h14];
  assign T399 = T79[5'h15:5'h15];
  assign T400 = T79[5'h16:5'h16];
  assign T401 = T79[5'h17:5'h17];
  assign T402 = T79[5'h18:5'h18];
  assign T403 = T79[5'h19:5'h19];
  assign T404 = T79[5'h1a:5'h1a];
  assign T405 = T79[5'h1b:5'h1b];
  assign T406 = T79[5'h1c:5'h1c];
  assign T407 = T79[5'h1d:5'h1d];
  assign T408 = T79[5'h1e:5'h1e];
  assign T409 = T79[5'h1f:5'h1f];
  assign T410 = T79[6'h20:6'h20];
  assign T411 = T79[6'h21:6'h21];
  assign T412 = T79[6'h22:6'h22];
  assign T413 = T79[6'h23:6'h23];
  assign T414 = T79[6'h24:6'h24];
  assign T415 = T79[6'h25:6'h25];
  assign T416 = T79[6'h26:6'h26];
  assign T417 = T79[6'h27:6'h27];
  assign T418 = T79[6'h28:6'h28];
  assign T419 = T79[6'h29:6'h29];
  assign T420 = T79[6'h2a:6'h2a];
  assign T421 = T79[6'h2b:6'h2b];
  assign T422 = T79[6'h2c:6'h2c];
  assign T423 = T79[6'h2d:6'h2d];
  assign T424 = T79[6'h2e:6'h2e];
  assign T425 = T79[6'h2f:6'h2f];
  assign T426 = T79[6'h30:6'h30];
  assign T427 = T79[6'h31:6'h31];
  assign T428 = T79[6'h32:6'h32];
  assign T429 = T79[6'h33:6'h33];
  assign T430 = T79[6'h34:6'h34];
  assign T431 = T79[6'h35:6'h35];
  assign T432 = T79[6'h36:6'h36];
  assign T433 = T79[6'h37:6'h37];
  assign T434 = T79[6'h38:6'h38];
  assign T435 = T79[6'h39:6'h39];
  assign T436 = T79[6'h3a:6'h3a];
  assign T437 = T79[6'h3b:6'h3b];
  assign T438 = T79[6'h3c:6'h3c];
  assign T439 = T79[6'h3d:6'h3d];
  assign T440 = T79[6'h3e:6'h3e];
  assign T441 = T79[6'h3f:6'h3f];
  assign T81 = T192 < T317;
  assign T82 = T94 & T83;
  assign T83 = cmdHi ? lhs_sign : T84;
  assign T84 = lhs_sign != rhs_sign;
  assign lhs_sign = lhsSigned & T85;
  assign T85 = T88 ? T87 : T86;
  assign T86 = io_req_bits_in1[5'h1f:5'h1f];
  assign T87 = io_req_bits_in1[6'h3f:6'h3f];
  assign T88 = 1'h1 == T89;
  assign T89 = io_req_bits_dw & 1'h1;
  assign lhsSigned = T90;
  assign T90 = T93 | T91;
  assign T91 = T92 == 4'h0;
  assign T92 = io_req_bits_fn & 4'h3;
  assign T93 = T61 | T17;
  assign T94 = cmdMul ^ 1'h1;
  assign T95 = isHi ? 3'h3 : 3'h5;
  assign T96 = T153 & T97;
  assign T97 = T99 | T98;
  assign T98 = count == 7'h7;
  assign T99 = T111 & T100;
  assign T100 = T101 == 64'h0;
  assign T101 = T107 & T102;
  assign T102 = ~ T103;
  assign T103 = T104[6'h3f:1'h0];
  assign T104 = $signed(65'h10000000000000000) >>> T105;
  assign T105 = T106[3'h5:1'h0];
  assign T106 = count * 4'h8;
  assign T107 = T108[6'h3f:1'h0];
  assign T108 = {T110, T109};
  assign T109 = remainder[6'h3f:1'h0];
  assign T110 = remainder[8'h81:7'h41];
  assign T111 = T113 & T112;
  assign T112 = isHi ^ 1'h1;
  assign T113 = T115 & T114;
  assign T114 = count != 7'h0;
  assign T115 = count != 7'h7;
  assign T116 = isHi ? 3'h3 : T117;
  assign T117 = neg_out ? 3'h4 : 3'h5;
  assign T118 = T162 & T119;
  assign T119 = count == 7'h40;
  assign T120 = T121 | io_kill;
  assign T121 = io_resp_ready & io_resp_valid;
  assign T122 = T123 ? 3'h1 : 3'h2;
  assign T123 = lhs_sign | T124;
  assign T124 = rhs_sign & T125;
  assign T125 = cmdMul ^ 1'h1;
  assign T442 = {66'h0, negated_remainder};
  assign T127 = state == 3'h4;
  assign T443 = {66'h0, T128};
  assign T128 = remainder[8'h80:7'h41];
  assign T129 = state == 3'h3;
  assign T130 = {T152, T131};
  assign T131 = {1'h0, T132};
  assign T132 = T133[6'h3f:1'h0];
  assign T133 = {T151, T134};
  assign T134 = T135[6'h3f:1'h0];
  assign T135 = T99 ? T147 : T136;
  assign T136 = T137;
  assign T137 = {T139, T138};
  assign T138 = T107[6'h3f:4'h8];
  assign T139 = T142 + T444;
  assign T444 = {T445, T140};
  assign T140 = T141;
  assign T141 = T108[8'h80:7'h40];
  assign T445 = T446 ? 8'hff : 8'h0;
  assign T446 = T140[7'h40:7'h40];
  assign T142 = $signed(T146) * $signed(T143);
  assign T143 = T144;
  assign T144 = {1'h0, T145};
  assign T145 = T107[3'h7:1'h0];
  assign T146 = divisor;
  assign T147 = T108 >> T148;
  assign T148 = T149[3'h5:1'h0];
  assign T149 = 11'h40 - T150;
  assign T150 = count * 4'h8;
  assign T151 = T136[8'h80:7'h40];
  assign T152 = T133 >> 7'h40;
  assign T153 = T154 & isMul;
  assign T154 = state == 3'h2;
  assign T447 = {1'h0, T155};
  assign T155 = {T159, T156};
  assign T156 = {T158, T157};
  assign T157 = less ^ 1'h1;
  assign T158 = remainder[6'h3f:1'h0];
  assign T159 = less ? T161 : T160;
  assign T160 = subtractor[6'h3f:1'h0];
  assign T161 = remainder[7'h7f:7'h40];
  assign T162 = T164 & T163;
  assign T163 = isMul ^ 1'h1;
  assign T164 = state == 3'h2;
  assign T448 = {3'h0, T165};
  assign T165 = T166 << T71;
  assign T166 = remainder[6'h3f:1'h0];
  assign T167 = T162 & T168;
  assign T168 = T171 & T169;
  assign T169 = T170 | T81;
  assign T170 = 6'h0 < T73;
  assign T171 = T172 & less;
  assign T172 = count == 7'h0;
  assign T449 = {66'h0, lhs_in};
  assign lhs_in = {T174, T173};
  assign T173 = io_req_bits_in1[5'h1f:1'h0];
  assign T174 = T177 ? T176 : T175;
  assign T175 = 32'h0 - T450;
  assign T450 = {31'h0, lhs_sign};
  assign T176 = io_req_bits_in1[6'h3f:6'h20];
  assign T177 = 1'h1 == T178;
  assign T178 = io_req_bits_dw & 1'h1;
  assign T179 = {T181, T180};
  assign T180 = remainder[5'h1f:1'h0];
  assign T181 = 32'h0 - T451;
  assign T451 = {31'h0, T182};
  assign T182 = remainder[5'h1f:5'h1f];
  assign T183 = 1'h0 == T184;
  assign T184 = req_dw & 1'h1;
  assign T185 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T186;
  assign T186 = state == 3'h5;
  assign io_req_ready = T187;
  assign T187 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T449;
    end else if(T167) begin
      remainder <= T448;
    end else if(T162) begin
      remainder <= T447;
    end else if(T153) begin
      remainder <= T130;
    end else if(T129) begin
      remainder <= T443;
    end else if(T127) begin
      remainder <= T442;
    end else if(T11) begin
      remainder <= T188;
    end
    if(T1) begin
      isMul <= cmdMul;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T122;
    end else if(T120) begin
      state <= 3'h0;
    end else if(T118) begin
      state <= T116;
    end else if(T96) begin
      state <= T95;
    end else if(T129) begin
      state <= T28;
    end else if(T127) begin
      state <= 3'h5;
    end else if(T20) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T82;
    end else if(T31) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= cmdHi;
    end
    if(T1) begin
      divisor <= T48;
    end else if(T45) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T167) begin
      count <= T191;
    end else if(T162) begin
      count <= T70;
    end else if(T153) begin
      count <= T69;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module Rocket(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_csr_req_ready,
    input  io_host_csr_req_valid,
    input  io_host_csr_req_bits_rw,
    input [11:0] io_host_csr_req_bits_addr,
    input [63:0] io_host_csr_req_bits_data,
    input  io_host_csr_resp_ready,
    output io_host_csr_resp_valid,
    output[63:0] io_host_csr_resp_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_csr,
    output io_imem_req_valid,
    output[39:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [39:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data_0,
    input  io_imem_resp_bits_mask,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input  io_imem_btb_resp_bits_mask,
    input  io_imem_btb_resp_bits_bridx,
    input [38:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output io_imem_btb_update_bits_prediction_bits_mask,
    output io_imem_btb_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_btb_update_bits_prediction_bits_target,
    output[5:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[38:0] io_imem_btb_update_bits_pc,
    output[38:0] io_imem_btb_update_bits_target,
    //output io_imem_btb_update_bits_taken
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isReturn,
    output[38:0] io_imem_btb_update_bits_br_pc,
    output io_imem_bht_update_valid,
    output io_imem_bht_update_bits_prediction_valid,
    output io_imem_bht_update_bits_prediction_bits_taken,
    output io_imem_bht_update_bits_prediction_bits_mask,
    output io_imem_bht_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_bht_update_bits_prediction_bits_target,
    output[5:0] io_imem_bht_update_bits_prediction_bits_entry,
    output[6:0] io_imem_bht_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
    output[38:0] io_imem_bht_update_bits_pc,
    output io_imem_bht_update_bits_taken,
    output io_imem_bht_update_bits_mispredict,
    output io_imem_ras_update_valid,
    output io_imem_ras_update_bits_isCall,
    output io_imem_ras_update_bits_isReturn,
    output[38:0] io_imem_ras_update_bits_returnAddr,
    output io_imem_ras_update_bits_prediction_valid,
    output io_imem_ras_update_bits_prediction_bits_taken,
    output io_imem_ras_update_bits_prediction_bits_mask,
    output io_imem_ras_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_ras_update_bits_prediction_bits_target,
    output[5:0] io_imem_ras_update_bits_prediction_bits_entry,
    output[6:0] io_imem_ras_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
    output io_imem_invalidate,
    input [39:0] io_imem_npc,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output[39:0] io_dmem_req_bits_addr,
    output[8:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_kill,
    output io_dmem_req_bits_phys,
    output[63:0] io_dmem_req_bits_data,
    input  io_dmem_resp_valid,
    input [39:0] io_dmem_resp_bits_addr,
    input [8:0] io_dmem_resp_bits_tag,
    input [4:0] io_dmem_resp_bits_cmd,
    input [2:0] io_dmem_resp_bits_typ,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_word_bypass,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [8:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    output io_dmem_invalidate_lr,
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_status_sd,
    output[30:0] io_ptw_status_zero2,
    output io_ptw_status_sd_rv32,
    output[8:0] io_ptw_status_zero1,
    output[4:0] io_ptw_status_vm,
    output io_ptw_status_mprv,
    output[1:0] io_ptw_status_xs,
    output[1:0] io_ptw_status_fs,
    output[1:0] io_ptw_status_prv3,
    output io_ptw_status_ie3,
    output[1:0] io_ptw_status_prv2,
    output io_ptw_status_ie2,
    output[1:0] io_ptw_status_prv1,
    output io_ptw_status_ie1,
    output[1:0] io_ptw_status_prv,
    output io_ptw_status_ie,
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    output io_fpu_valid,
    //input  io_fpu_fcsr_rdy
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    //input [4:0] io_fpu_dec_cmd
    //input  io_fpu_dec_ldst
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    //input  io_fpu_dec_swap12
    //input  io_fpu_dec_swap23
    //input  io_fpu_dec_single
    //input  io_fpu_dec_fromint
    //input  io_fpu_dec_toint
    //input  io_fpu_dec_fastpipe
    //input  io_fpu_dec_fma
    //input  io_fpu_dec_div
    //input  io_fpu_dec_sqrt
    //input  io_fpu_dec_round
    //input  io_fpu_dec_wflags
    //input  io_fpu_sboard_set
    //input  io_fpu_sboard_clr
    //input [4:0] io_fpu_sboard_clra
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input [39:0] io_rocc_mem_req_bits_addr,
    input [8:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_kill,
    input  io_rocc_mem_req_bits_phys,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[39:0] io_rocc_mem_resp_bits_addr
    //output[8:0] io_rocc_mem_resp_bits_tag
    //output[4:0] io_rocc_mem_resp_bits_cmd
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_word_bypass
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[8:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_invalidate_lr,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [25:0] io_rocc_imem_acquire_bits_addr_block,
    input [1:0] io_rocc_imem_acquire_bits_client_xact_id,
    input [1:0] io_rocc_imem_acquire_bits_addr_beat,
    input  io_rocc_imem_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_imem_acquire_bits_a_type,
    input [16:0] io_rocc_imem_acquire_bits_union,
    input [127:0] io_rocc_imem_acquire_bits_data,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_addr_beat
    //output[1:0] io_rocc_imem_grant_bits_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_manager_xact_id
    //output io_rocc_imem_grant_bits_is_builtin_type
    //output[3:0] io_rocc_imem_grant_bits_g_type
    //output[127:0] io_rocc_imem_grant_bits_data
    //output io_rocc_dmem_0_acquire_ready
    input  io_rocc_dmem_0_acquire_valid,
    input [25:0] io_rocc_dmem_0_acquire_bits_addr_block,
    input [1:0] io_rocc_dmem_0_acquire_bits_client_xact_id,
    input [1:0] io_rocc_dmem_0_acquire_bits_addr_beat,
    input  io_rocc_dmem_0_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_dmem_0_acquire_bits_a_type,
    input [16:0] io_rocc_dmem_0_acquire_bits_union,
    input [127:0] io_rocc_dmem_0_acquire_bits_data,
    input  io_rocc_dmem_0_grant_ready,
    //output io_rocc_dmem_0_grant_valid
    //output[1:0] io_rocc_dmem_0_grant_bits_addr_beat
    //output[1:0] io_rocc_dmem_0_grant_bits_client_xact_id
    //output[3:0] io_rocc_dmem_0_grant_bits_manager_xact_id
    //output io_rocc_dmem_0_grant_bits_is_builtin_type
    //output[3:0] io_rocc_dmem_0_grant_bits_g_type
    //output[127:0] io_rocc_dmem_0_grant_bits_data
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [26:0] io_rocc_iptw_req_bits_addr,
    input [1:0] io_rocc_iptw_req_bits_prv,
    input  io_rocc_iptw_req_bits_store,
    input  io_rocc_iptw_req_bits_fetch,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[19:0] io_rocc_iptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_iptw_resp_bits_pte_reserved_for_software
    //output io_rocc_iptw_resp_bits_pte_d
    //output io_rocc_iptw_resp_bits_pte_r
    //output[3:0] io_rocc_iptw_resp_bits_pte_typ
    //output io_rocc_iptw_resp_bits_pte_v
    //output io_rocc_iptw_status_sd
    //output[30:0] io_rocc_iptw_status_zero2
    //output io_rocc_iptw_status_sd_rv32
    //output[8:0] io_rocc_iptw_status_zero1
    //output[4:0] io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_mprv
    //output[1:0] io_rocc_iptw_status_xs
    //output[1:0] io_rocc_iptw_status_fs
    //output[1:0] io_rocc_iptw_status_prv3
    //output io_rocc_iptw_status_ie3
    //output[1:0] io_rocc_iptw_status_prv2
    //output io_rocc_iptw_status_ie2
    //output[1:0] io_rocc_iptw_status_prv1
    //output io_rocc_iptw_status_ie1
    //output[1:0] io_rocc_iptw_status_prv
    //output io_rocc_iptw_status_ie
    //output io_rocc_iptw_invalidate
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [26:0] io_rocc_dptw_req_bits_addr,
    input [1:0] io_rocc_dptw_req_bits_prv,
    input  io_rocc_dptw_req_bits_store,
    input  io_rocc_dptw_req_bits_fetch,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[19:0] io_rocc_dptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_dptw_resp_bits_pte_reserved_for_software
    //output io_rocc_dptw_resp_bits_pte_d
    //output io_rocc_dptw_resp_bits_pte_r
    //output[3:0] io_rocc_dptw_resp_bits_pte_typ
    //output io_rocc_dptw_resp_bits_pte_v
    //output io_rocc_dptw_status_sd
    //output[30:0] io_rocc_dptw_status_zero2
    //output io_rocc_dptw_status_sd_rv32
    //output[8:0] io_rocc_dptw_status_zero1
    //output[4:0] io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_mprv
    //output[1:0] io_rocc_dptw_status_xs
    //output[1:0] io_rocc_dptw_status_fs
    //output[1:0] io_rocc_dptw_status_prv3
    //output io_rocc_dptw_status_ie3
    //output[1:0] io_rocc_dptw_status_prv2
    //output io_rocc_dptw_status_ie2
    //output[1:0] io_rocc_dptw_status_prv1
    //output io_rocc_dptw_status_ie1
    //output[1:0] io_rocc_dptw_status_prv
    //output io_rocc_dptw_status_ie
    //output io_rocc_dptw_invalidate
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [26:0] io_rocc_pptw_req_bits_addr,
    input [1:0] io_rocc_pptw_req_bits_prv,
    input  io_rocc_pptw_req_bits_store,
    input  io_rocc_pptw_req_bits_fetch,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[19:0] io_rocc_pptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_pptw_resp_bits_pte_reserved_for_software
    //output io_rocc_pptw_resp_bits_pte_d
    //output io_rocc_pptw_resp_bits_pte_r
    //output[3:0] io_rocc_pptw_resp_bits_pte_typ
    //output io_rocc_pptw_resp_bits_pte_v
    //output io_rocc_pptw_status_sd
    //output[30:0] io_rocc_pptw_status_zero2
    //output io_rocc_pptw_status_sd_rv32
    //output[8:0] io_rocc_pptw_status_zero1
    //output[4:0] io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_mprv
    //output[1:0] io_rocc_pptw_status_xs
    //output[1:0] io_rocc_pptw_status_fs
    //output[1:0] io_rocc_pptw_status_prv3
    //output io_rocc_pptw_status_ie3
    //output[1:0] io_rocc_pptw_status_prv2
    //output io_rocc_pptw_status_ie2
    //output[1:0] io_rocc_pptw_status_prv1
    //output io_rocc_pptw_status_ie1
    //output[1:0] io_rocc_pptw_status_prv
    //output io_rocc_pptw_status_ie
    //output io_rocc_pptw_invalidate
    output io_rocc_exception
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  wire ctrl_killd;
  wire T7;
  wire T8;
  wire ctrl_stalld;
  wire T9;
  wire id_do_fence;
  wire T10;
  wire id_csr_en;
  wire[2:0] id_ctrl_csr;
  wire[2:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[31:0] T14;
  wire T15;
  wire[31:0] T16;
  wire T17;
  wire[31:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire id_ctrl_rocc;
  wire id_ctrl_mem;
  wire T22;
  wire T23;
  wire[31:0] T24;
  wire T25;
  wire T26;
  wire[31:0] T27;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire T31;
  wire T32;
  wire[31:0] T33;
  wire T34;
  wire T35;
  wire[31:0] T36;
  wire T37;
  wire[31:0] T38;
  reg  id_reg_fence;
  wire T916;
  wire T39;
  wire T40;
  wire id_fence_next;
  wire T41;
  wire id_amo_rl;
  wire id_ctrl_amo;
  wire T42;
  wire[31:0] T43;
  wire id_ctrl_fence;
  wire T44;
  wire[31:0] T45;
  wire T46;
  wire id_ctrl_fence_i;
  wire T47;
  wire[31:0] T48;
  wire T49;
  wire id_amo_aq;
  wire id_mem_busy;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire id_sboard_hazard;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[4:0] T59;
  wire[4:0] T60;
  wire[4:0] id_waddr;
  wire T61;
  wire[31:0] T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire[31:0] T65;
  wire[4:0] ll_waddr;
  wire[4:0] T66;
  wire[4:0] dmem_resp_waddr;
  wire[8:0] T67;
  wire T68;
  wire dmem_resp_xpu;
  wire T69;
  wire T70;
  wire dmem_resp_replay;
  wire ll_wen;
  wire T71;
  wire T72;
  reg [31:0] R73;
  wire[31:0] T917;
  wire[31:0] T74;
  wire[31:0] T75;
  wire[31:0] T76;
  wire[31:0] T77;
  wire[31:0] T78;
  wire[4:0] wb_waddr;
  wire T79;
  wire wb_wen;
  reg  wb_ctrl_wxd;
  wire T80;
  reg  mem_ctrl_wxd;
  wire T81;
  reg  ex_ctrl_wxd;
  wire T82;
  wire id_ctrl_wxd;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire T87;
  wire[31:0] T88;
  wire T89;
  wire T90;
  wire[31:0] T91;
  wire T92;
  wire T93;
  wire[31:0] T94;
  wire T95;
  wire T96;
  wire[31:0] T97;
  wire T98;
  wire T99;
  wire[31:0] T100;
  wire T101;
  wire[31:0] T102;
  wire T103;
  wire wb_valid;
  wire T104;
  wire T105;
  wire T106;
  wire replay_wb;
  wire T107;
  wire T108;
  wire T109;
  reg  wb_ctrl_rocc;
  wire T110;
  reg  mem_ctrl_rocc;
  wire T111;
  reg  ex_ctrl_rocc;
  wire T112;
  wire replay_wb_common;
  wire T113;
  reg  wb_reg_replay;
  wire T114;
  wire T115;
  wire take_pc_wb;
  wire T116;
  wire T117;
  wire wb_xcpt;
  reg  wb_reg_xcpt;
  wire T118;
  wire T119;
  wire mem_xcpt;
  wire T120;
  wire T121;
  reg  mem_ctrl_mem;
  wire T122;
  reg  ex_ctrl_mem;
  wire T123;
  reg  mem_reg_valid;
  wire T124;
  wire ctrl_killx;
  wire T125;
  reg  ex_reg_valid;
  wire T126;
  wire T127;
  wire replay_ex;
  wire T128;
  wire replay_ex_load_use;
  reg  ex_reg_load_use;
  wire T129;
  wire id_load_use;
  wire T130;
  wire T131;
  wire data_hazard_mem;
  wire T132;
  wire T133;
  wire T134;
  wire[4:0] mem_waddr;
  wire T135;
  wire T136;
  wire T137;
  wire[4:0] id_raddr_1;
  wire T138;
  wire T139;
  wire id_ctrl_rxs2;
  wire T140;
  wire T141;
  wire[31:0] T142;
  wire T143;
  wire T144;
  wire[31:0] T145;
  wire T146;
  wire[31:0] T147;
  wire T148;
  wire T149;
  wire[4:0] id_raddr_0;
  wire T150;
  wire T151;
  wire id_ctrl_rxs1;
  wire T152;
  wire T153;
  wire[31:0] T154;
  wire T155;
  wire T156;
  wire[31:0] T157;
  wire T158;
  wire T159;
  wire[31:0] T160;
  wire T161;
  wire[31:0] T162;
  wire wb_dcache_miss;
  wire T163;
  reg  wb_ctrl_mem;
  wire T164;
  wire replay_ex_structural;
  wire T165;
  wire T166;
  reg  ex_ctrl_div;
  wire T167;
  wire id_ctrl_div;
  wire T168;
  wire[31:0] T169;
  wire T170;
  wire T171;
  wire take_pc;
  wire take_pc_mem;
  wire T172;
  wire T173;
  wire mem_npc_misaligned;
  wire[39:0] mem_npc;
  wire[39:0] T174;
  wire[39:0] T175;
  wire[39:0] mem_br_target;
  wire[39:0] T918;
  wire[21:0] T176;
  wire[21:0] T177;
  wire[21:0] T178;
  wire[21:0] T179;
  wire[11:0] T180;
  wire[4:0] T181;
  wire[3:0] T182;
  wire[6:0] T183;
  wire[5:0] T184;
  wire T185;
  wire T186;
  wire[9:0] T187;
  wire[8:0] T188;
  wire[7:0] T189;
  wire[7:0] T190;
  wire T191;
  wire T192;
  reg  mem_ctrl_jal;
  wire T193;
  reg  ex_ctrl_jal;
  wire T194;
  wire id_ctrl_jal;
  wire[21:0] T919;
  wire[14:0] T195;
  wire[14:0] T196;
  wire[11:0] T197;
  wire[4:0] T198;
  wire[3:0] T199;
  wire[6:0] T200;
  wire[5:0] T201;
  wire T202;
  wire T203;
  wire[2:0] T204;
  wire[1:0] T205;
  wire T206;
  wire T207;
  wire[6:0] T920;
  wire T921;
  wire T208;
  wire mem_br_taken;
  reg [63:0] bypass_mux_1;
  wire[63:0] T209;
  reg  mem_ctrl_branch;
  wire T210;
  reg  ex_ctrl_branch;
  wire T211;
  wire id_ctrl_branch;
  wire T212;
  wire[31:0] T213;
  wire[17:0] T922;
  wire T923;
  wire[39:0] T214;
  reg [39:0] mem_reg_pc;
  wire[39:0] T215;
  reg [39:0] ex_reg_pc;
  wire[39:0] T216;
  wire[39:0] T217;
  wire[39:0] T218;
  wire[38:0] T219;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire[1:0] T225;
  wire T226;
  wire T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire T230;
  wire[25:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  reg  mem_ctrl_jalr;
  wire T236;
  reg  ex_ctrl_jalr;
  wire T237;
  wire id_ctrl_jalr;
  wire T238;
  wire[31:0] T239;
  wire want_take_pc_mem;
  wire T240;
  reg  mem_reg_flush_pipe;
  wire T241;
  reg  ex_reg_flush_pipe;
  wire T242;
  wire T243;
  wire id_csr_flush;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[11:0] T248;
  wire[11:0] id_csr_addr;
  wire T249;
  wire T250;
  wire id_csr_ren;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire id_system_insn;
  wire mem_misprediction;
  wire T255;
  wire T256;
  wire T257;
  wire mem_wrong_npc;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  reg  mem_reg_xcpt;
  wire T272;
  wire ex_xcpt;
  wire T273;
  reg  ex_ctrl_fp;
  wire T274;
  wire id_ctrl_fp;
  wire T275;
  reg  ex_reg_xcpt;
  wire T276;
  wire id_xcpt;
  wire id_illegal_insn;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire id_ctrl_legal;
  wire T285;
  wire T286;
  wire[31:0] T287;
  wire T288;
  wire T289;
  wire[31:0] T290;
  wire T291;
  wire T292;
  wire[31:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[31:0] T298;
  wire T299;
  wire T300;
  wire T301;
  wire[31:0] T302;
  wire T303;
  wire T304;
  wire T305;
  wire[31:0] T306;
  wire T307;
  wire T308;
  wire[31:0] T309;
  wire T310;
  wire T311;
  wire[31:0] T312;
  wire T313;
  wire T314;
  wire[31:0] T315;
  wire T316;
  wire T317;
  wire[31:0] T318;
  wire T319;
  wire T320;
  wire T321;
  wire[31:0] T322;
  wire T323;
  wire T324;
  wire[31:0] T325;
  wire T326;
  wire T327;
  wire[31:0] T328;
  wire T329;
  wire T330;
  wire[31:0] T331;
  wire T332;
  wire T333;
  wire[31:0] T334;
  wire T335;
  wire T336;
  wire[31:0] T337;
  wire T338;
  wire T339;
  wire[31:0] T340;
  wire T341;
  wire T342;
  wire[31:0] T343;
  wire T344;
  wire T345;
  wire[31:0] T346;
  wire T347;
  wire T348;
  wire[31:0] T349;
  wire T350;
  wire T351;
  wire[31:0] T352;
  wire T353;
  wire T354;
  wire[31:0] T355;
  wire T356;
  wire T357;
  wire T358;
  reg  ex_reg_xcpt_interrupt;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  reg  mem_reg_xcpt_interrupt;
  wire T363;
  wire T364;
  wire replay_mem;
  wire fpu_kill_mem;
  wire T365;
  reg  mem_ctrl_fp;
  wire T366;
  wire T367;
  reg  mem_reg_replay;
  wire T368;
  wire T369;
  wire dcache_kill_mem;
  wire T370;
  reg  wb_reg_valid;
  wire T371;
  wire ctrl_killm;
  wire T372;
  wire killm_common;
  wire T373;
  wire T374;
  wire T375;
  wire wb_set_sboard;
  wire T376;
  reg  wb_ctrl_div;
  wire T377;
  reg  mem_ctrl_div;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire[4:0] T387;
  wire[4:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[4:0] T394;
  wire[4:0] T395;
  wire T396;
  wire T397;
  wire id_wb_hazard;
  wire T398;
  wire fp_data_hazard_wb;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire[4:0] id_raddr3;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  reg  wb_ctrl_wfd;
  wire T410;
  reg  mem_ctrl_wfd;
  wire T411;
  reg  ex_ctrl_wfd;
  wire T412;
  wire id_ctrl_wfd;
  wire T413;
  wire data_hazard_wb;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire id_mem_hazard;
  wire T423;
  wire fp_data_hazard_mem;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire mem_cannot_bypass;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  reg  mem_mem_cmd_bh;
  wire T440;
  wire ex_slow_bypass;
  wire T441;
  wire T442;
  reg [2:0] ex_ctrl_mem_type;
  wire[2:0] T443;
  wire[2:0] id_ctrl_mem_type;
  wire[2:0] T444;
  wire[1:0] T445;
  wire T446;
  wire[31:0] T447;
  wire T448;
  wire[31:0] T449;
  wire T450;
  wire[31:0] T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  reg [4:0] ex_ctrl_mem_cmd;
  wire[4:0] T458;
  wire[4:0] id_ctrl_mem_cmd;
  wire[4:0] T459;
  wire[3:0] T460;
  wire[2:0] T461;
  wire[1:0] T462;
  wire T463;
  wire T464;
  wire[31:0] T465;
  wire T466;
  wire T467;
  wire[31:0] T468;
  wire T469;
  wire[31:0] T470;
  wire T471;
  wire T472;
  wire[31:0] T473;
  wire T474;
  wire[31:0] T475;
  wire T476;
  wire T477;
  wire[31:0] T478;
  wire T479;
  wire T480;
  wire[31:0] T481;
  wire T482;
  wire[31:0] T483;
  wire T484;
  reg [2:0] mem_ctrl_csr;
  wire[2:0] T485;
  reg [2:0] ex_ctrl_csr;
  wire[2:0] T486;
  wire[2:0] T487;
  wire[2:0] id_csr;
  wire id_ex_hazard;
  wire T488;
  wire fp_data_hazard_ex;
  wire T489;
  wire T490;
  wire T491;
  wire[4:0] ex_waddr;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire ex_cannot_bypass;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire data_hazard_ex;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire[31:0] T519;
  wire[63:0] T520;
  reg [63:0] R521;
  reg [63:0] R522;
  wire[63:0] ex_rs_1;
  wire[63:0] T523;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T524;
  wire[1:0] T525;
  wire[1:0] T526;
  wire[1:0] T527;
  wire[1:0] T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire[1:0] T538;
  wire[63:0] id_rs_1;
  wire[63:0] T539;
  wire[63:0] T540;
  reg [63:0] T541 [30:0];
  wire[63:0] T542;
  wire T543;
  wire T544;
  wire[4:0] T545;
  wire T546;
  wire T547;
  wire[4:0] rf_waddr;
  wire rf_wen;
  wire[4:0] T548;
  wire[4:0] T549;
  wire[63:0] rf_wdata;
  wire[63:0] T550;
  wire[63:0] T551;
  reg [63:0] bypass_mux_2;
  wire[63:0] T552;
  wire[63:0] T553;
  wire[63:0] mem_int_wdata;
  wire[63:0] T554;
  wire[63:0] T555;
  wire[63:0] T924;
  wire[23:0] T925;
  wire T926;
  wire T556;
  wire T557;
  reg [2:0] wb_ctrl_csr;
  wire[2:0] T558;
  wire[63:0] ll_wdata;
  wire T559;
  wire dmem_resp_valid;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T571;
  wire[61:0] T572;
  wire[63:0] T573;
  wire[63:0] T574;
  wire T575;
  wire[1:0] T576;
  wire[63:0] T577;
  wire T578;
  wire T579;
  reg  ex_reg_rs_bypass_1;
  wire T580;
  wire[4:0] T581;
  wire[4:0] T582;
  wire[63:0] T583;
  reg [63:0] R584;
  reg [63:0] R585;
  wire[63:0] ex_rs_0;
  wire[63:0] T586;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire[1:0] T590;
  wire[1:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[1:0] T597;
  wire[63:0] id_rs_0;
  wire[63:0] T598;
  wire[63:0] T599;
  wire[4:0] T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T611;
  wire[61:0] T612;
  wire[63:0] T613;
  wire[63:0] T614;
  wire T615;
  wire[1:0] T616;
  wire[63:0] T617;
  wire T618;
  wire T619;
  reg  ex_reg_rs_bypass_0;
  wire T620;
  wire[4:0] T621;
  wire[4:0] T622;
  wire T623;
  wire[63:0] T624;
  wire[4:0] T625;
  wire[4:0] T626;
  wire[39:0] T627;
  reg [39:0] wb_reg_pc;
  wire[39:0] T628;
  wire T629;
  wire[32:0] T630;
  wire[32:0] T631;
  wire T632;
  wire[1127:0] T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  reg  R638;
  wire T639;
  reg  ex_ctrl_alu_dw;
  wire T640;
  wire id_ctrl_alu_dw;
  wire T641;
  wire T642;
  wire[31:0] T643;
  wire T644;
  wire[31:0] T645;
  reg [3:0] ex_ctrl_alu_fn;
  wire[3:0] T646;
  wire[3:0] id_ctrl_alu_fn;
  wire[3:0] T647;
  wire[2:0] T648;
  wire[1:0] T649;
  wire T650;
  wire T651;
  wire[31:0] T652;
  wire T653;
  wire T654;
  wire[31:0] T655;
  wire T656;
  wire[31:0] T657;
  wire T658;
  wire T659;
  wire[31:0] T660;
  wire T661;
  wire T662;
  wire[31:0] T663;
  wire T664;
  wire T665;
  wire[31:0] T666;
  wire T667;
  wire T668;
  wire[31:0] T669;
  wire T670;
  wire[31:0] T671;
  wire T672;
  wire T673;
  wire[31:0] T674;
  wire T675;
  wire T676;
  wire[31:0] T677;
  wire T678;
  wire T679;
  wire[31:0] T680;
  wire T681;
  wire[31:0] T682;
  wire T683;
  wire T684;
  wire[31:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire[31:0] T689;
  wire T690;
  wire[63:0] T691;
  wire[63:0] ex_op1;
  wire[63:0] T927;
  wire[39:0] T692;
  wire[39:0] T693;
  wire T694;
  reg [1:0] ex_ctrl_sel_alu1;
  wire[1:0] T695;
  wire[1:0] id_ctrl_sel_alu1;
  wire[1:0] T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire[31:0] T701;
  wire T702;
  wire T703;
  wire[31:0] T704;
  wire[23:0] T928;
  wire T929;
  wire[63:0] T705;
  wire T706;
  wire[63:0] T707;
  wire[63:0] ex_op2;
  wire[63:0] T930;
  wire[31:0] T708;
  wire[31:0] T931;
  wire[3:0] T709;
  wire T710;
  reg [1:0] ex_ctrl_sel_alu2;
  wire[1:0] T711;
  wire[1:0] id_ctrl_sel_alu2;
  wire[1:0] T712;
  wire T713;
  wire T714;
  wire[31:0] T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire[31:0] T720;
  wire T721;
  wire[31:0] T722;
  wire T723;
  wire T724;
  wire[31:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[31:0] T729;
  wire[27:0] T932;
  wire T933;
  wire[31:0] ex_imm;
  wire[31:0] T730;
  wire[11:0] T731;
  wire[4:0] T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  reg [2:0] ex_ctrl_sel_imm;
  wire[2:0] T738;
  wire[2:0] id_ctrl_sel_imm;
  wire[2:0] T739;
  wire[1:0] T740;
  wire T741;
  wire T742;
  wire[31:0] T743;
  wire T744;
  wire[31:0] T745;
  wire T746;
  wire T747;
  wire[31:0] T748;
  wire T749;
  wire T750;
  wire[31:0] T751;
  wire T752;
  wire T753;
  wire[31:0] T754;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[3:0] T759;
  wire[3:0] T760;
  wire[3:0] T761;
  wire[3:0] T762;
  wire[3:0] T763;
  wire T764;
  wire[3:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire[6:0] T770;
  wire[5:0] T771;
  wire[5:0] T772;
  wire T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire T791;
  wire[19:0] T792;
  wire[18:0] T793;
  wire[7:0] T794;
  wire[7:0] T795;
  wire[7:0] T796;
  wire[7:0] T934;
  wire T797;
  wire T798;
  wire T799;
  wire[10:0] T800;
  wire[10:0] T935;
  wire[10:0] T801;
  wire[10:0] T802;
  wire T803;
  wire T804;
  wire[31:0] T936;
  wire T937;
  wire[63:0] T805;
  wire T806;
  reg [63:0] wb_reg_cause;
  wire[63:0] T807;
  wire[63:0] mem_cause;
  wire[63:0] T938;
  wire[2:0] T808;
  wire[2:0] T809;
  wire[2:0] T810;
  wire[2:0] T811;
  reg [63:0] mem_reg_cause;
  wire[63:0] T812;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T813;
  wire[63:0] id_cause;
  wire[63:0] T939;
  wire[1:0] T814;
  wire[2:0] T815;
  wire[11:0] T816;
  wire T817;
  wire T818;
  wire T819;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T820;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T821;
  wire T822;
  wire T823;
  wire T824;
  reg  ex_ctrl_rxs2;
  wire T825;
  wire T826;
  wire[6:0] T827;
  wire[4:0] T828;
  wire T829;
  wire T830;
  wire T831;
  wire[4:0] T832;
  wire[4:0] T833;
  wire[6:0] T834;
  wire wb_rocc_val;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire dmem_resp_fpu;
  wire T840;
  wire[63:0] T841;
  wire T842;
  wire[8:0] T940;
  wire[5:0] T843;
  wire[39:0] T844;
  wire[39:0] T845;
  wire[38:0] T846;
  wire T847;
  wire T848;
  wire T849;
  wire[1:0] T850;
  wire T851;
  wire[1:0] T852;
  wire T853;
  wire T854;
  wire[25:0] T855;
  wire[25:0] T856;
  wire T857;
  wire[25:0] T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  reg  wb_ctrl_fence_i;
  wire T865;
  reg  mem_ctrl_fence_i;
  wire T866;
  reg  ex_ctrl_fence_i;
  wire T867;
  wire[38:0] T941;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire[38:0] T942;
  wire T875;
  wire T876;
  wire T877;
  wire[38:0] T943;
  wire T878;
  wire T879;
  wire[4:0] T880;
  wire[4:0] T881;
  wire T882;
  wire[38:0] T944;
  wire[38:0] T945;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T883;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T884;
  wire T885;
  wire T886;
  reg  ex_reg_btb_hit;
  wire T887;
  reg [6:0] mem_reg_btb_resp_bht_history;
  wire[6:0] T888;
  reg [6:0] ex_reg_btb_resp_bht_history;
  wire[6:0] T889;
  reg [5:0] mem_reg_btb_resp_entry;
  wire[5:0] T890;
  reg [5:0] ex_reg_btb_resp_entry;
  wire[5:0] T891;
  reg [38:0] mem_reg_btb_resp_target;
  wire[38:0] T892;
  reg [38:0] ex_reg_btb_resp_target;
  wire[38:0] T893;
  reg  mem_reg_btb_resp_bridx;
  wire T894;
  reg  ex_reg_btb_resp_bridx;
  wire T895;
  reg  mem_reg_btb_resp_mask;
  wire T896;
  reg  ex_reg_btb_resp_mask;
  wire T897;
  reg  mem_reg_btb_resp_taken;
  wire T898;
  reg  ex_reg_btb_resp_taken;
  wire T899;
  reg  mem_reg_btb_hit;
  wire T900;
  wire T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire T911;
  wire[39:0] T912;
  wire[39:0] T913;
  wire[39:0] T914;
  wire T915;
  wire csr_io_host_csr_req_ready;
  wire csr_io_host_csr_resp_valid;
  wire[63:0] csr_io_host_csr_resp_bits;
  wire csr_io_host_ipi_req_valid;
  wire csr_io_host_ipi_req_bits;
  wire csr_io_host_ipi_rep_ready;
  wire csr_io_host_debug_stats_csr;
  wire[63:0] csr_io_rw_rdata;
  wire csr_io_csr_replay;
  wire csr_io_csr_stall;
  wire csr_io_csr_xcpt;
  wire csr_io_eret;
  wire csr_io_status_sd;
  wire[30:0] csr_io_status_zero2;
  wire csr_io_status_sd_rv32;
  wire[8:0] csr_io_status_zero1;
  wire[4:0] csr_io_status_vm;
  wire csr_io_status_mprv;
  wire[1:0] csr_io_status_xs;
  wire[1:0] csr_io_status_fs;
  wire[1:0] csr_io_status_prv3;
  wire csr_io_status_ie3;
  wire[1:0] csr_io_status_prv2;
  wire csr_io_status_ie2;
  wire[1:0] csr_io_status_prv1;
  wire csr_io_status_ie1;
  wire[1:0] csr_io_status_prv;
  wire csr_io_status_ie;
  wire[31:0] csr_io_ptbr;
  wire[39:0] csr_io_evec;
  wire csr_io_fatc;
  wire[63:0] csr_io_time;
  wire[2:0] csr_io_fcsr_rm;
  wire csr_io_interrupt;
  wire[63:0] csr_io_interrupt_cause;
  wire[63:0] alu_io_out;
  wire[63:0] alu_io_adder_out;
  wire div_io_req_ready;
  wire div_io_resp_valid;
  wire[63:0] div_io_resp_bits_data;
  wire[4:0] div_io_resp_bits_tag;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    id_reg_fence = {1{$random}};
    R73 = {1{$random}};
    wb_ctrl_wxd = {1{$random}};
    mem_ctrl_wxd = {1{$random}};
    ex_ctrl_wxd = {1{$random}};
    wb_ctrl_rocc = {1{$random}};
    mem_ctrl_rocc = {1{$random}};
    ex_ctrl_rocc = {1{$random}};
    wb_reg_replay = {1{$random}};
    wb_reg_xcpt = {1{$random}};
    mem_ctrl_mem = {1{$random}};
    ex_ctrl_mem = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    ex_reg_load_use = {1{$random}};
    wb_ctrl_mem = {1{$random}};
    ex_ctrl_div = {1{$random}};
    mem_ctrl_jal = {1{$random}};
    ex_ctrl_jal = {1{$random}};
    bypass_mux_1 = {2{$random}};
    mem_ctrl_branch = {1{$random}};
    ex_ctrl_branch = {1{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    mem_ctrl_jalr = {1{$random}};
    ex_ctrl_jalr = {1{$random}};
    mem_reg_flush_pipe = {1{$random}};
    ex_reg_flush_pipe = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_ctrl_fp = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    mem_ctrl_fp = {1{$random}};
    mem_reg_replay = {1{$random}};
    wb_reg_valid = {1{$random}};
    wb_ctrl_div = {1{$random}};
    mem_ctrl_div = {1{$random}};
    wb_ctrl_wfd = {1{$random}};
    mem_ctrl_wfd = {1{$random}};
    ex_ctrl_wfd = {1{$random}};
    mem_mem_cmd_bh = {1{$random}};
    ex_ctrl_mem_type = {1{$random}};
    ex_ctrl_mem_cmd = {1{$random}};
    mem_ctrl_csr = {1{$random}};
    ex_ctrl_csr = {1{$random}};
    R521 = {2{$random}};
    R522 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T541[initvar] = {2{$random}};
    bypass_mux_2 = {2{$random}};
    wb_ctrl_csr = {1{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R584 = {2{$random}};
    R585 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    R638 = {1{$random}};
    ex_ctrl_alu_dw = {1{$random}};
    ex_ctrl_alu_fn = {1{$random}};
    ex_ctrl_sel_alu1 = {1{$random}};
    ex_ctrl_sel_alu2 = {1{$random}};
    ex_ctrl_sel_imm = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
    ex_ctrl_rxs2 = {1{$random}};
    wb_ctrl_fence_i = {1{$random}};
    mem_ctrl_fence_i = {1{$random}};
    ex_ctrl_fence_i = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_history = {1{$random}};
    ex_reg_btb_resp_bht_history = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_bridx = {1{$random}};
    ex_reg_btb_resp_bridx = {1{$random}};
    mem_reg_btb_resp_mask = {1{$random}};
    ex_reg_btb_resp_mask = {1{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_ie = {1{$random}};
//  assign io_rocc_pptw_status_prv = {1{$random}};
//  assign io_rocc_pptw_status_ie1 = {1{$random}};
//  assign io_rocc_pptw_status_prv1 = {1{$random}};
//  assign io_rocc_pptw_status_ie2 = {1{$random}};
//  assign io_rocc_pptw_status_prv2 = {1{$random}};
//  assign io_rocc_pptw_status_ie3 = {1{$random}};
//  assign io_rocc_pptw_status_prv3 = {1{$random}};
//  assign io_rocc_pptw_status_fs = {1{$random}};
//  assign io_rocc_pptw_status_xs = {1{$random}};
//  assign io_rocc_pptw_status_mprv = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_zero1 = {1{$random}};
//  assign io_rocc_pptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_pptw_status_zero2 = {1{$random}};
//  assign io_rocc_pptw_status_sd = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_ie = {1{$random}};
//  assign io_rocc_dptw_status_prv = {1{$random}};
//  assign io_rocc_dptw_status_ie1 = {1{$random}};
//  assign io_rocc_dptw_status_prv1 = {1{$random}};
//  assign io_rocc_dptw_status_ie2 = {1{$random}};
//  assign io_rocc_dptw_status_prv2 = {1{$random}};
//  assign io_rocc_dptw_status_ie3 = {1{$random}};
//  assign io_rocc_dptw_status_prv3 = {1{$random}};
//  assign io_rocc_dptw_status_fs = {1{$random}};
//  assign io_rocc_dptw_status_xs = {1{$random}};
//  assign io_rocc_dptw_status_mprv = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_zero1 = {1{$random}};
//  assign io_rocc_dptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_dptw_status_zero2 = {1{$random}};
//  assign io_rocc_dptw_status_sd = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_ie = {1{$random}};
//  assign io_rocc_iptw_status_prv = {1{$random}};
//  assign io_rocc_iptw_status_ie1 = {1{$random}};
//  assign io_rocc_iptw_status_prv1 = {1{$random}};
//  assign io_rocc_iptw_status_ie2 = {1{$random}};
//  assign io_rocc_iptw_status_prv2 = {1{$random}};
//  assign io_rocc_iptw_status_ie3 = {1{$random}};
//  assign io_rocc_iptw_status_prv3 = {1{$random}};
//  assign io_rocc_iptw_status_fs = {1{$random}};
//  assign io_rocc_iptw_status_xs = {1{$random}};
//  assign io_rocc_iptw_status_mprv = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_zero1 = {1{$random}};
//  assign io_rocc_iptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_iptw_status_zero2 = {1{$random}};
//  assign io_rocc_iptw_status_sd = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_data = {4{$random}};
//  assign io_rocc_dmem_0_grant_bits_g_type = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_dmem_0_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_dmem_0_grant_valid = {1{$random}};
//  assign io_rocc_dmem_0_acquire_ready = {1{$random}};
//  assign io_rocc_imem_grant_bits_data = {4{$random}};
//  assign io_rocc_imem_grant_bits_g_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_imem_grant_valid = {1{$random}};
//  assign io_rocc_imem_acquire_ready = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_data_word_bypass = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
//  assign io_imem_btb_update_bits_taken = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T517 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T516 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data_0 : ex_reg_inst;
  assign T5 = T6 | csr_io_interrupt;
  assign T6 = ctrl_killd ^ 1'h1;
  assign ctrl_killd = T7;
  assign T7 = T8 | csr_io_interrupt;
  assign T8 = T514 | ctrl_stalld;
  assign ctrl_stalld = T9 | csr_io_csr_stall;
  assign T9 = T51 | id_do_fence;
  assign id_do_fence = id_mem_busy & T10;
  assign T10 = T19 | id_csr_en;
  assign id_csr_en = id_ctrl_csr != 3'h0;
  assign id_ctrl_csr = T11;
  assign T11 = {T17, T12};
  assign T12 = {T15, T13};
  assign T13 = T14 == 32'h1050;
  assign T14 = io_imem_resp_bits_data_0 & 32'h1050;
  assign T15 = T16 == 32'h2050;
  assign T16 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T17 = T18 == 32'h50;
  assign T18 = io_imem_resp_bits_data_0 & 32'h3050;
  assign T19 = T46 | T20;
  assign T20 = id_reg_fence & T21;
  assign T21 = id_ctrl_mem | id_ctrl_rocc;
  assign id_ctrl_rocc = 1'h0;
  assign id_ctrl_mem = T22;
  assign T22 = T25 | T23;
  assign T23 = T24 == 32'h1000202f;
  assign T24 = io_imem_resp_bits_data_0 & 32'hf9f0607f;
  assign T25 = T28 | T26;
  assign T26 = T27 == 32'h800202f;
  assign T27 = io_imem_resp_bits_data_0 & 32'he800607f;
  assign T28 = T31 | T29;
  assign T29 = T30 == 32'h202f;
  assign T30 = io_imem_resp_bits_data_0 & 32'h1800607f;
  assign T31 = T34 | T32;
  assign T32 = T33 == 32'h3;
  assign T33 = io_imem_resp_bits_data_0 & 32'h107f;
  assign T34 = T37 | T35;
  assign T35 = T36 == 32'h3;
  assign T36 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T37 = T38 == 32'h3;
  assign T38 = io_imem_resp_bits_data_0 & 32'h405f;
  assign T916 = reset ? 1'h0 : T39;
  assign T39 = id_fence_next | T40;
  assign T40 = id_reg_fence & id_mem_busy;
  assign id_fence_next = id_ctrl_fence | T41;
  assign T41 = id_ctrl_amo & id_amo_rl;
  assign id_amo_rl = io_imem_resp_bits_data_0[5'h19:5'h19];
  assign id_ctrl_amo = T42;
  assign T42 = T43 == 32'h2008;
  assign T43 = io_imem_resp_bits_data_0 & 32'h6048;
  assign id_ctrl_fence = T44;
  assign T44 = T45 == 32'h8;
  assign T45 = io_imem_resp_bits_data_0 & 32'h3058;
  assign T46 = T49 | id_ctrl_fence_i;
  assign id_ctrl_fence_i = T47;
  assign T47 = T48 == 32'h1008;
  assign T48 = io_imem_resp_bits_data_0 & 32'h3058;
  assign T49 = id_ctrl_amo & id_amo_aq;
  assign id_amo_aq = io_imem_resp_bits_data_0[5'h1a:5'h1a];
  assign id_mem_busy = T50 | io_dmem_req_valid;
  assign T50 = io_dmem_ordered ^ 1'h1;
  assign T51 = T54 | T52;
  assign T52 = id_ctrl_mem & T53;
  assign T53 = io_dmem_req_ready ^ 1'h1;
  assign T54 = T397 | id_sboard_hazard;
  assign id_sboard_hazard = T382 | T55;
  assign T55 = T380 & T56;
  assign T56 = T61 & T57;
  assign T57 = T58 - 1'h1;
  assign T58 = 1'h1 << T59;
  assign T59 = T60 + 5'h1;
  assign T60 = id_waddr - id_waddr;
  assign id_waddr = io_imem_resp_bits_data_0[4'hb:3'h7];
  assign T61 = T62 >> id_waddr;
  assign T62 = R73 & T63;
  assign T63 = ~ T64;
  assign T64 = ll_wen ? T65 : 32'h0;
  assign T65 = 1'h1 << ll_waddr;
  assign ll_waddr = T66;
  assign T66 = T68 ? dmem_resp_waddr : div_io_resp_bits_tag;
  assign dmem_resp_waddr = T67[3'h5:1'h1];
  assign T67 = io_dmem_resp_bits_tag;
  assign T68 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_xpu = T69 ^ 1'h1;
  assign T69 = T70;
  assign T70 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign ll_wen = T71;
  assign T71 = T68 ? 1'h1 : T72;
  assign T72 = T634 & div_io_resp_valid;
  assign T917 = reset ? 32'h0 : T74;
  assign T74 = T379 ? T76 : T75;
  assign T75 = ll_wen ? T62 : R73;
  assign T76 = T62 | T77;
  assign T77 = T79 ? T78 : 32'h0;
  assign T78 = 1'h1 << wb_waddr;
  assign wb_waddr = wb_reg_inst[4'hb:3'h7];
  assign T79 = wb_set_sboard & wb_wen;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign T80 = T517 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign T81 = T516 ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign T82 = T103 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign id_ctrl_wxd = T83;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h0;
  assign T85 = io_imem_resp_bits_data_0 & 32'h28;
  assign T86 = T89 | T87;
  assign T87 = T88 == 32'h2010;
  assign T88 = io_imem_resp_bits_data_0 & 32'h2010;
  assign T89 = T92 | T90;
  assign T90 = T91 == 32'h2008;
  assign T91 = io_imem_resp_bits_data_0 & 32'h2008;
  assign T92 = T95 | T93;
  assign T93 = T94 == 32'h1010;
  assign T94 = io_imem_resp_bits_data_0 & 32'h1010;
  assign T95 = T98 | T96;
  assign T96 = T97 == 32'h48;
  assign T97 = io_imem_resp_bits_data_0 & 32'h48;
  assign T98 = T101 | T99;
  assign T99 = T100 == 32'h10;
  assign T100 = io_imem_resp_bits_data_0 & 32'h50;
  assign T101 = T102 == 32'h4;
  assign T102 = io_imem_resp_bits_data_0 & 32'hc;
  assign T103 = ctrl_killd ^ 1'h1;
  assign wb_valid = T105 & T104;
  assign T104 = csr_io_csr_xcpt ^ 1'h1;
  assign T105 = wb_reg_valid & T106;
  assign T106 = replay_wb ^ 1'h1;
  assign replay_wb = replay_wb_common | T107;
  assign T107 = T109 & T108;
  assign T108 = io_rocc_cmd_ready ^ 1'h1;
  assign T109 = wb_reg_valid & wb_ctrl_rocc;
  assign T110 = T517 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign T111 = T516 ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign T112 = T103 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign replay_wb_common = T113 | csr_io_csr_replay;
  assign T113 = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T114 = replay_mem & T115;
  assign T115 = take_pc_wb ^ 1'h1;
  assign take_pc_wb = T116;
  assign T116 = T117 | csr_io_eret;
  assign T117 = replay_wb | wb_xcpt;
  assign wb_xcpt = wb_reg_xcpt | csr_io_csr_xcpt;
  assign T118 = mem_xcpt & T119;
  assign T119 = take_pc_wb ^ 1'h1;
  assign mem_xcpt = T260 | T120;
  assign T120 = T121 & io_dmem_xcpt_pf_ld;
  assign T121 = mem_reg_valid & mem_ctrl_mem;
  assign T122 = T516 ? ex_ctrl_mem : mem_ctrl_mem;
  assign T123 = T103 ? id_ctrl_mem : ex_ctrl_mem;
  assign T124 = ctrl_killx ^ 1'h1;
  assign ctrl_killx = T127 | T125;
  assign T125 = ex_reg_valid ^ 1'h1;
  assign T126 = ctrl_killd ^ 1'h1;
  assign T127 = take_pc | replay_ex;
  assign replay_ex = ex_reg_valid & T128;
  assign T128 = replay_ex_structural | replay_ex_load_use;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T129 = T103 ? id_load_use : ex_reg_load_use;
  assign id_load_use = T130;
  assign T130 = T131 & mem_ctrl_mem;
  assign T131 = mem_reg_valid & data_hazard_mem;
  assign data_hazard_mem = mem_ctrl_wxd & T132;
  assign T132 = T135 | T133;
  assign T133 = T380 & T134;
  assign T134 = id_waddr == mem_waddr;
  assign mem_waddr = mem_reg_inst[4'hb:3'h7];
  assign T135 = T148 | T136;
  assign T136 = T138 & T137;
  assign T137 = id_raddr_1 == mem_waddr;
  assign id_raddr_1 = io_imem_resp_bits_data_0[5'h18:5'h14];
  assign T138 = id_ctrl_rxs2 & T139;
  assign T139 = id_raddr_1 != 5'h0;
  assign id_ctrl_rxs2 = T140;
  assign T140 = T143 | T141;
  assign T141 = T142 == 32'h20;
  assign T142 = io_imem_resp_bits_data_0 & 32'h34;
  assign T143 = T146 | T144;
  assign T144 = T145 == 32'h20;
  assign T145 = io_imem_resp_bits_data_0 & 32'h64;
  assign T146 = T147 == 32'h20;
  assign T147 = io_imem_resp_bits_data_0 & 32'h70;
  assign T148 = T150 & T149;
  assign T149 = id_raddr_0 == mem_waddr;
  assign id_raddr_0 = io_imem_resp_bits_data_0[5'h13:4'hf];
  assign T150 = id_ctrl_rxs1 & T151;
  assign T151 = id_raddr_0 != 5'h0;
  assign id_ctrl_rxs1 = T152;
  assign T152 = T155 | T153;
  assign T153 = T154 == 32'h2000;
  assign T154 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T155 = T158 | T156;
  assign T156 = T157 == 32'h0;
  assign T157 = io_imem_resp_bits_data_0 & 32'h18;
  assign T158 = T161 | T159;
  assign T159 = T160 == 32'h0;
  assign T160 = io_imem_resp_bits_data_0 & 32'h44;
  assign T161 = T162 == 32'h0;
  assign T162 = io_imem_resp_bits_data_0 & 32'h4004;
  assign wb_dcache_miss = wb_ctrl_mem & T163;
  assign T163 = io_dmem_resp_valid ^ 1'h1;
  assign T164 = T517 ? mem_ctrl_mem : wb_ctrl_mem;
  assign replay_ex_structural = T170 | T165;
  assign T165 = ex_ctrl_div & T166;
  assign T166 = div_io_req_ready ^ 1'h1;
  assign T167 = T103 ? id_ctrl_div : ex_ctrl_div;
  assign id_ctrl_div = T168;
  assign T168 = T169 == 32'h2000030;
  assign T169 = io_imem_resp_bits_data_0 & 32'h2000074;
  assign T170 = ex_ctrl_mem & T171;
  assign T171 = io_dmem_req_ready ^ 1'h1;
  assign take_pc = take_pc_wb | take_pc_mem;
  assign take_pc_mem = T172;
  assign T172 = want_take_pc_mem & T173;
  assign T173 = mem_npc_misaligned ^ 1'h1;
  assign mem_npc_misaligned = mem_npc[1'h1:1'h1];
  assign mem_npc = T174;
  assign T174 = T175 & 40'hfffffffffe;
  assign T175 = mem_ctrl_jalr ? T217 : mem_br_target;
  assign mem_br_target = T214 + T918;
  assign T918 = {T922, T176};
  assign T176 = T208 ? T919 : T177;
  assign T177 = mem_ctrl_jal ? T178 : 22'h4;
  assign T178 = T179;
  assign T179 = {T187, T180};
  assign T180 = {T183, T181};
  assign T181 = {T182, 1'h0};
  assign T182 = mem_reg_inst[5'h18:5'h15];
  assign T183 = {T185, T184};
  assign T184 = mem_reg_inst[5'h1e:5'h19];
  assign T185 = T186;
  assign T186 = mem_reg_inst[5'h14:5'h14];
  assign T187 = {T191, T188};
  assign T188 = {T191, T189};
  assign T189 = T190;
  assign T190 = mem_reg_inst[5'h13:4'hc];
  assign T191 = T192;
  assign T192 = mem_reg_inst[5'h1f:5'h1f];
  assign T193 = T516 ? ex_ctrl_jal : mem_ctrl_jal;
  assign T194 = T103 ? id_ctrl_jal : ex_ctrl_jal;
  assign id_ctrl_jal = T96;
  assign T919 = {T920, T195};
  assign T195 = T196;
  assign T196 = {T204, T197};
  assign T197 = {T200, T198};
  assign T198 = {T199, 1'h0};
  assign T199 = mem_reg_inst[4'hb:4'h8];
  assign T200 = {T202, T201};
  assign T201 = mem_reg_inst[5'h1e:5'h19];
  assign T202 = T203;
  assign T203 = mem_reg_inst[3'h7:3'h7];
  assign T204 = {T206, T205};
  assign T205 = {T206, T206};
  assign T206 = T207;
  assign T207 = mem_reg_inst[5'h1f:5'h1f];
  assign T920 = T921 ? 7'h7f : 7'h0;
  assign T921 = T195[4'he:4'he];
  assign T208 = mem_ctrl_branch & mem_br_taken;
  assign mem_br_taken = bypass_mux_1[1'h0:1'h0];
  assign T209 = T516 ? alu_io_out : bypass_mux_1;
  assign T210 = T516 ? ex_ctrl_branch : mem_ctrl_branch;
  assign T211 = T103 ? id_ctrl_branch : ex_ctrl_branch;
  assign id_ctrl_branch = T212;
  assign T212 = T213 == 32'h40;
  assign T213 = io_imem_resp_bits_data_0 & 32'h54;
  assign T922 = T923 ? 18'h3ffff : 18'h0;
  assign T923 = T176[5'h15:5'h15];
  assign T214 = mem_reg_pc;
  assign T215 = T516 ? ex_reg_pc : mem_reg_pc;
  assign T216 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T217 = T218;
  assign T218 = {T220, T219};
  assign T219 = bypass_mux_1[6'h26:1'h0];
  assign T220 = T233 ? T232 : T221;
  assign T221 = T226 ? T224 : T222;
  assign T222 = T223[1'h0:1'h0];
  assign T223 = bypass_mux_1[6'h27:6'h26];
  assign T224 = T225 == 2'h3;
  assign T225 = T223;
  assign T226 = T230 | T227;
  assign T227 = T228 == 26'h3fffffe;
  assign T228 = T229;
  assign T229 = bypass_mux_1 >> 6'h26;
  assign T230 = T231 == 26'h3ffffff;
  assign T231 = T229;
  assign T232 = T223 != 2'h0;
  assign T233 = T235 | T234;
  assign T234 = T229 == 26'h1;
  assign T235 = T229 == 26'h0;
  assign T236 = T516 ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign T237 = T103 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign id_ctrl_jalr = T238;
  assign T238 = T239 == 32'h4;
  assign T239 = io_imem_resp_bits_data_0 & 32'h1c;
  assign want_take_pc_mem = mem_reg_valid & T240;
  assign T240 = mem_misprediction | mem_reg_flush_pipe;
  assign T241 = T516 ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign T242 = T103 ? T243 : ex_reg_flush_pipe;
  assign T243 = id_ctrl_fence_i | id_csr_flush;
  assign id_csr_flush = id_system_insn | T244;
  assign T244 = T249 & T245;
  assign T245 = T246 ^ 1'h1;
  assign T246 = T247;
  assign T247 = T248 == 12'h40;
  assign T248 = id_csr_addr & 12'h8c4;
  assign id_csr_addr = io_imem_resp_bits_data_0[5'h1f:5'h14];
  assign T249 = id_csr_en & T250;
  assign T250 = id_csr_ren ^ 1'h1;
  assign id_csr_ren = T252 & T251;
  assign T251 = id_raddr_0 == 5'h0;
  assign T252 = T254 | T253;
  assign T253 = id_ctrl_csr == 3'h3;
  assign T254 = id_ctrl_csr == 3'h2;
  assign id_system_insn = id_ctrl_csr == 3'h4;
  assign mem_misprediction = T257 & T255;
  assign T255 = T256 | mem_ctrl_jal;
  assign T256 = mem_ctrl_branch | mem_ctrl_jalr;
  assign T257 = mem_wrong_npc & mem_reg_valid;
  assign mem_wrong_npc = T259 | T258;
  assign T258 = ex_reg_valid ^ 1'h1;
  assign T259 = mem_npc != ex_reg_pc;
  assign T260 = T263 | T261;
  assign T261 = T262 & io_dmem_xcpt_pf_st;
  assign T262 = mem_reg_valid & mem_ctrl_mem;
  assign T263 = T266 | T264;
  assign T264 = T265 & io_dmem_xcpt_ma_ld;
  assign T265 = mem_reg_valid & mem_ctrl_mem;
  assign T266 = T269 | T267;
  assign T267 = T268 & io_dmem_xcpt_ma_st;
  assign T268 = mem_reg_valid & mem_ctrl_mem;
  assign T269 = T271 | T270;
  assign T270 = want_take_pc_mem & mem_npc_misaligned;
  assign T271 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T272 = T362 & ex_xcpt;
  assign ex_xcpt = T275 | T273;
  assign T273 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign T274 = T103 ? id_ctrl_fp : ex_ctrl_fp;
  assign id_ctrl_fp = 1'h0;
  assign T275 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T276 = T358 & id_xcpt;
  assign id_xcpt = T357 | id_illegal_insn;
  assign id_illegal_insn = T280 | T277;
  assign T277 = id_ctrl_rocc & T278;
  assign T278 = T279 ^ 1'h1;
  assign T279 = csr_io_status_xs != 2'h0;
  assign T280 = T284 | T281;
  assign T281 = id_ctrl_fp & T282;
  assign T282 = T283 ^ 1'h1;
  assign T283 = csr_io_status_fs != 2'h0;
  assign T284 = id_ctrl_legal ^ 1'h1;
  assign id_ctrl_legal = T285;
  assign T285 = T288 | T286;
  assign T286 = T287 == 32'h33;
  assign T287 = io_imem_resp_bits_data_0 & 32'hfc007077;
  assign T288 = T291 | T289;
  assign T289 = T290 == 32'h4063;
  assign T290 = io_imem_resp_bits_data_0 & 32'h407f;
  assign T291 = T294 | T292;
  assign T292 = T293 == 32'h1063;
  assign T293 = io_imem_resp_bits_data_0 & 32'h306f;
  assign T294 = T296 | T295;
  assign T295 = io_imem_resp_bits_data_0 == 32'h30500073;
  assign T296 = T299 | T297;
  assign T297 = T298 == 32'h10100073;
  assign T298 = io_imem_resp_bits_data_0 & 32'hfff07fff;
  assign T299 = T300 | T23;
  assign T300 = T303 | T301;
  assign T301 = T302 == 32'h10000073;
  assign T302 = io_imem_resp_bits_data_0 & 32'hffdfffff;
  assign T303 = T304 | T26;
  assign T304 = T307 | T305;
  assign T305 = T306 == 32'h2004033;
  assign T306 = io_imem_resp_bits_data_0 & 32'hfe004077;
  assign T307 = T310 | T308;
  assign T308 = T309 == 32'h5033;
  assign T309 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T310 = T313 | T311;
  assign T311 = T312 == 32'h501b;
  assign T312 = io_imem_resp_bits_data_0 & 32'hbe00705f;
  assign T313 = T316 | T314;
  assign T314 = T315 == 32'h5013;
  assign T315 = io_imem_resp_bits_data_0 & 32'hbc00707f;
  assign T316 = T319 | T317;
  assign T317 = T318 == 32'h2073;
  assign T318 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T319 = T320 | T29;
  assign T320 = T323 | T321;
  assign T321 = T322 == 32'h2013;
  assign T322 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T323 = T326 | T324;
  assign T324 = T325 == 32'h101b;
  assign T325 = io_imem_resp_bits_data_0 & 32'hfe00305f;
  assign T326 = T329 | T327;
  assign T327 = T328 == 32'h1013;
  assign T328 = io_imem_resp_bits_data_0 & 32'hfc00305f;
  assign T329 = T332 | T330;
  assign T330 = T331 == 32'h73;
  assign T331 = io_imem_resp_bits_data_0 & 32'hffefffff;
  assign T332 = T335 | T333;
  assign T333 = T334 == 32'h6f;
  assign T334 = io_imem_resp_bits_data_0 & 32'h7f;
  assign T335 = T338 | T336;
  assign T336 = T337 == 32'h63;
  assign T337 = io_imem_resp_bits_data_0 & 32'h707b;
  assign T338 = T341 | T339;
  assign T339 = T340 == 32'h33;
  assign T340 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T341 = T344 | T342;
  assign T342 = T343 == 32'h33;
  assign T343 = io_imem_resp_bits_data_0 & 32'hfc00007f;
  assign T344 = T347 | T345;
  assign T345 = T346 == 32'h17;
  assign T346 = io_imem_resp_bits_data_0 & 32'h5f;
  assign T347 = T350 | T348;
  assign T348 = T349 == 32'h13;
  assign T349 = io_imem_resp_bits_data_0 & 32'h7077;
  assign T350 = T353 | T351;
  assign T351 = T352 == 32'hf;
  assign T352 = io_imem_resp_bits_data_0 & 32'h607f;
  assign T353 = T356 | T354;
  assign T354 = T355 == 32'h3;
  assign T355 = io_imem_resp_bits_data_0 & 32'h106f;
  assign T356 = T37 | T35;
  assign T357 = csr_io_interrupt | io_imem_resp_bits_xcpt_if;
  assign T358 = ctrl_killd ^ 1'h1;
  assign T359 = T360 & io_imem_resp_valid;
  assign T360 = csr_io_interrupt & T361;
  assign T361 = take_pc ^ 1'h1;
  assign T362 = ctrl_killx ^ 1'h1;
  assign T363 = T364 & ex_reg_xcpt_interrupt;
  assign T364 = take_pc ^ 1'h1;
  assign replay_mem = T367 | fpu_kill_mem;
  assign fpu_kill_mem = T365 & io_fpu_nack_mem;
  assign T365 = mem_reg_valid & mem_ctrl_fp;
  assign T366 = T516 ? ex_ctrl_fp : mem_ctrl_fp;
  assign T367 = dcache_kill_mem | mem_reg_replay;
  assign T368 = T369 & replay_ex;
  assign T369 = take_pc ^ 1'h1;
  assign dcache_kill_mem = T370 & io_dmem_replay_next_valid;
  assign T370 = mem_reg_valid & mem_ctrl_wxd;
  assign T371 = ctrl_killm ^ 1'h1;
  assign ctrl_killm = T372 | fpu_kill_mem;
  assign T372 = killm_common | mem_xcpt;
  assign killm_common = T374 | T373;
  assign T373 = mem_reg_valid ^ 1'h1;
  assign T374 = T375 | mem_reg_xcpt;
  assign T375 = dcache_kill_mem | take_pc_wb;
  assign wb_set_sboard = T376 | wb_ctrl_rocc;
  assign T376 = wb_ctrl_div | wb_dcache_miss;
  assign T377 = T517 ? mem_ctrl_div : wb_ctrl_div;
  assign T378 = T516 ? ex_ctrl_div : mem_ctrl_div;
  assign T379 = ll_wen | T79;
  assign T380 = id_ctrl_wxd & T381;
  assign T381 = id_waddr != 5'h0;
  assign T382 = T390 | T383;
  assign T383 = T138 & T384;
  assign T384 = T389 & T385;
  assign T385 = T386 - 1'h1;
  assign T386 = 1'h1 << T387;
  assign T387 = T388 + 5'h1;
  assign T388 = id_raddr_1 - id_raddr_1;
  assign T389 = T62 >> id_raddr_1;
  assign T390 = T150 & T391;
  assign T391 = T396 & T392;
  assign T392 = T393 - 1'h1;
  assign T393 = 1'h1 << T394;
  assign T394 = T395 + 5'h1;
  assign T395 = id_raddr_0 - id_raddr_0;
  assign T396 = T62 >> id_raddr_0;
  assign T397 = T422 | id_wb_hazard;
  assign id_wb_hazard = wb_reg_valid & T398;
  assign T398 = T413 | fp_data_hazard_wb;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T399;
  assign T399 = T402 | T400;
  assign T400 = io_fpu_dec_wen & T401;
  assign T401 = id_waddr == wb_waddr;
  assign T402 = T405 | T403;
  assign T403 = io_fpu_dec_ren3 & T404;
  assign T404 = id_raddr3 == wb_waddr;
  assign id_raddr3 = io_imem_resp_bits_data_0[5'h1f:5'h1b];
  assign T405 = T408 | T406;
  assign T406 = io_fpu_dec_ren2 & T407;
  assign T407 = id_raddr_1 == wb_waddr;
  assign T408 = io_fpu_dec_ren1 & T409;
  assign T409 = id_raddr_0 == wb_waddr;
  assign T410 = T517 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign T411 = T516 ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign T412 = T103 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign id_ctrl_wfd = 1'h0;
  assign T413 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_ctrl_wxd & T414;
  assign T414 = T417 | T415;
  assign T415 = T380 & T416;
  assign T416 = id_waddr == wb_waddr;
  assign T417 = T420 | T418;
  assign T418 = T138 & T419;
  assign T419 = id_raddr_1 == wb_waddr;
  assign T420 = T150 & T421;
  assign T421 = id_raddr_0 == wb_waddr;
  assign T422 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = mem_reg_valid & T423;
  assign T423 = T435 | fp_data_hazard_mem;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T424;
  assign T424 = T427 | T425;
  assign T425 = io_fpu_dec_wen & T426;
  assign T426 = id_waddr == mem_waddr;
  assign T427 = T430 | T428;
  assign T428 = io_fpu_dec_ren3 & T429;
  assign T429 = id_raddr3 == mem_waddr;
  assign T430 = T433 | T431;
  assign T431 = io_fpu_dec_ren2 & T432;
  assign T432 = id_raddr_1 == mem_waddr;
  assign T433 = io_fpu_dec_ren1 & T434;
  assign T434 = id_raddr_0 == mem_waddr;
  assign T435 = data_hazard_mem & mem_cannot_bypass;
  assign mem_cannot_bypass = T436 | mem_ctrl_rocc;
  assign T436 = T437 | mem_ctrl_fp;
  assign T437 = T438 | mem_ctrl_div;
  assign T438 = T484 | T439;
  assign T439 = mem_ctrl_mem & mem_mem_cmd_bh;
  assign T440 = T516 ? ex_slow_bypass : mem_mem_cmd_bh;
  assign ex_slow_bypass = T457 | T441;
  assign T441 = T452 | T442;
  assign T442 = 3'h5 == ex_ctrl_mem_type;
  assign T443 = T103 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign id_ctrl_mem_type = T444;
  assign T444 = {T450, T445};
  assign T445 = {T448, T446};
  assign T446 = T447 == 32'h1000;
  assign T447 = io_imem_resp_bits_data_0 & 32'h1000;
  assign T448 = T449 == 32'h2000;
  assign T449 = io_imem_resp_bits_data_0 & 32'h2000;
  assign T450 = T451 == 32'h4000;
  assign T451 = io_imem_resp_bits_data_0 & 32'h4000;
  assign T452 = T454 | T453;
  assign T453 = 3'h1 == ex_ctrl_mem_type;
  assign T454 = T456 | T455;
  assign T455 = 3'h4 == ex_ctrl_mem_type;
  assign T456 = 3'h0 == ex_ctrl_mem_type;
  assign T457 = ex_ctrl_mem_cmd == 5'h7;
  assign T458 = T103 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign id_ctrl_mem_cmd = T459;
  assign T459 = {1'h0, T460};
  assign T460 = {T482, T461};
  assign T461 = {T476, T462};
  assign T462 = {T471, T463};
  assign T463 = T466 | T464;
  assign T464 = T465 == 32'h20000020;
  assign T465 = io_imem_resp_bits_data_0 & 32'h20000020;
  assign T466 = T469 | T467;
  assign T467 = T468 == 32'h18000020;
  assign T468 = io_imem_resp_bits_data_0 & 32'h18000020;
  assign T469 = T470 == 32'h20;
  assign T470 = io_imem_resp_bits_data_0 & 32'h28;
  assign T471 = T474 | T472;
  assign T472 = T473 == 32'h40000008;
  assign T473 = io_imem_resp_bits_data_0 & 32'h40000008;
  assign T474 = T475 == 32'h10000008;
  assign T475 = io_imem_resp_bits_data_0 & 32'h10000008;
  assign T476 = T479 | T477;
  assign T477 = T478 == 32'h80000008;
  assign T478 = io_imem_resp_bits_data_0 & 32'h80000008;
  assign T479 = T480 | T474;
  assign T480 = T481 == 32'h8000008;
  assign T481 = io_imem_resp_bits_data_0 & 32'h8000008;
  assign T482 = T483 == 32'h8;
  assign T483 = io_imem_resp_bits_data_0 & 32'h18000008;
  assign T484 = mem_ctrl_csr != 3'h0;
  assign T485 = T516 ? ex_ctrl_csr : mem_ctrl_csr;
  assign T486 = T103 ? id_csr : T487;
  assign T487 = T103 ? id_ctrl_csr : ex_ctrl_csr;
  assign id_csr = id_csr_ren ? 3'h5 : id_ctrl_csr;
  assign id_ex_hazard = ex_reg_valid & T488;
  assign T488 = T500 | fp_data_hazard_ex;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T489;
  assign T489 = T492 | T490;
  assign T490 = io_fpu_dec_wen & T491;
  assign T491 = id_waddr == ex_waddr;
  assign ex_waddr = ex_reg_inst[4'hb:3'h7];
  assign T492 = T495 | T493;
  assign T493 = io_fpu_dec_ren3 & T494;
  assign T494 = id_raddr3 == ex_waddr;
  assign T495 = T498 | T496;
  assign T496 = io_fpu_dec_ren2 & T497;
  assign T497 = id_raddr_1 == ex_waddr;
  assign T498 = io_fpu_dec_ren1 & T499;
  assign T499 = id_raddr_0 == ex_waddr;
  assign T500 = data_hazard_ex & ex_cannot_bypass;
  assign ex_cannot_bypass = T501 | ex_ctrl_rocc;
  assign T501 = T502 | ex_ctrl_fp;
  assign T502 = T503 | ex_ctrl_div;
  assign T503 = T504 | ex_ctrl_mem;
  assign T504 = T505 | ex_ctrl_jalr;
  assign T505 = ex_ctrl_csr != 3'h0;
  assign data_hazard_ex = ex_ctrl_wxd & T506;
  assign T506 = T509 | T507;
  assign T507 = T380 & T508;
  assign T508 = id_waddr == ex_waddr;
  assign T509 = T512 | T510;
  assign T510 = T138 & T511;
  assign T511 = id_raddr_1 == ex_waddr;
  assign T512 = T150 & T513;
  assign T513 = id_raddr_0 == ex_waddr;
  assign T514 = T515 | take_pc;
  assign T515 = io_imem_resp_valid ^ 1'h1;
  assign T516 = ex_reg_valid | ex_reg_xcpt_interrupt;
  assign T517 = T518 | mem_reg_xcpt_interrupt;
  assign T518 = mem_reg_valid | mem_reg_replay;
  assign T519 = wb_reg_inst;
  assign T520 = R521;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T573 : T523;
  assign T523 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T524 = T562 ? T538 : T525;
  assign T525 = T103 ? T526 : ex_reg_rs_lsb_1;
  assign T526 = T537 ? 2'h0 : T527;
  assign T527 = T534 ? 2'h1 : T528;
  assign T528 = T529 ? 2'h2 : 2'h3;
  assign T529 = T531 & T530;
  assign T530 = mem_waddr == id_raddr_1;
  assign T531 = T533 & T532;
  assign T532 = mem_ctrl_mem ^ 1'h1;
  assign T533 = mem_reg_valid & mem_ctrl_wxd;
  assign T534 = T536 & T535;
  assign T535 = ex_waddr == id_raddr_1;
  assign T536 = ex_reg_valid & ex_ctrl_wxd;
  assign T537 = 5'h0 == id_raddr_1;
  assign T538 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T539;
  assign T539 = T560 ? rf_wdata : T540;
  assign T540 = T541[T549];
  assign T543 = T546 & T544;
  assign T544 = T545 < 5'h1f;
  assign T545 = T548[3'h4:1'h0];
  assign T546 = rf_wen & T547;
  assign T547 = rf_waddr != 5'h0;
  assign rf_waddr = ll_wen ? ll_waddr : wb_waddr;
  assign rf_wen = wb_wen | ll_wen;
  assign T548 = ~ rf_waddr;
  assign T549 = ~ id_raddr_1;
  assign rf_wdata = T559 ? io_dmem_resp_bits_data : T550;
  assign T550 = ll_wen ? ll_wdata : T551;
  assign T551 = T557 ? csr_io_rw_rdata : bypass_mux_2;
  assign T552 = T517 ? T553 : bypass_mux_2;
  assign T553 = T556 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = T554;
  assign T554 = mem_ctrl_jalr ? T924 : T555;
  assign T555 = bypass_mux_1;
  assign T924 = {T925, mem_br_target};
  assign T925 = T926 ? 24'hffffff : 24'h0;
  assign T926 = mem_br_target[6'h27:6'h27];
  assign T556 = mem_ctrl_fp & mem_ctrl_wxd;
  assign T557 = wb_ctrl_csr != 3'h0;
  assign T558 = T517 ? mem_ctrl_csr : wb_ctrl_csr;
  assign ll_wdata = div_io_resp_bits_data;
  assign T559 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T560 = T546 & T561;
  assign T561 = rf_waddr == id_raddr_1;
  assign T562 = T103 & T563;
  assign T563 = id_ctrl_rxs2 & T564;
  assign T564 = T565 ^ 1'h1;
  assign T565 = T569 | T566;
  assign T566 = T568 & T567;
  assign T567 = mem_waddr == id_raddr_1;
  assign T568 = mem_reg_valid & mem_ctrl_wxd;
  assign T569 = T570 | T529;
  assign T570 = T537 | T534;
  assign T571 = T562 ? T572 : ex_reg_rs_msb_1;
  assign T572 = id_rs_1 >> 2'h2;
  assign T573 = T579 ? T577 : T574;
  assign T574 = T575 ? bypass_mux_1 : 64'h0;
  assign T575 = T576[1'h0:1'h0];
  assign T576 = ex_reg_rs_lsb_1;
  assign T577 = T578 ? io_dmem_resp_bits_data_word_bypass : bypass_mux_2;
  assign T578 = T576[1'h0:1'h0];
  assign T579 = T576[1'h1:1'h1];
  assign T580 = T103 ? T565 : ex_reg_rs_bypass_1;
  assign T581 = T582;
  assign T582 = wb_reg_inst[5'h18:5'h14];
  assign T583 = R584;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T613 : T586;
  assign T586 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T587 = T603 ? T597 : T588;
  assign T588 = T103 ? T589 : ex_reg_rs_lsb_0;
  assign T589 = T596 ? 2'h0 : T590;
  assign T590 = T594 ? 2'h1 : T591;
  assign T591 = T592 ? 2'h2 : 2'h3;
  assign T592 = T531 & T593;
  assign T593 = mem_waddr == id_raddr_0;
  assign T594 = T536 & T595;
  assign T595 = ex_waddr == id_raddr_0;
  assign T596 = 5'h0 == id_raddr_0;
  assign T597 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T598;
  assign T598 = T601 ? rf_wdata : T599;
  assign T599 = T541[T600];
  assign T600 = ~ id_raddr_0;
  assign T601 = T546 & T602;
  assign T602 = rf_waddr == id_raddr_0;
  assign T603 = T103 & T604;
  assign T604 = id_ctrl_rxs1 & T605;
  assign T605 = T606 ^ 1'h1;
  assign T606 = T609 | T607;
  assign T607 = T568 & T608;
  assign T608 = mem_waddr == id_raddr_0;
  assign T609 = T610 | T592;
  assign T610 = T596 | T594;
  assign T611 = T603 ? T612 : ex_reg_rs_msb_0;
  assign T612 = id_rs_0 >> 2'h2;
  assign T613 = T619 ? T617 : T614;
  assign T614 = T615 ? bypass_mux_1 : 64'h0;
  assign T615 = T616[1'h0:1'h0];
  assign T616 = ex_reg_rs_lsb_0;
  assign T617 = T618 ? io_dmem_resp_bits_data_word_bypass : bypass_mux_2;
  assign T618 = T616[1'h0:1'h0];
  assign T619 = T616[1'h1:1'h1];
  assign T620 = T103 ? T606 : ex_reg_rs_bypass_0;
  assign T621 = T622;
  assign T622 = wb_reg_inst[5'h13:4'hf];
  assign T623 = rf_wen;
  assign T624 = rf_wdata;
  assign T625 = T626;
  assign T626 = rf_wen ? rf_waddr : 5'h0;
  assign T627 = wb_reg_pc;
  assign T628 = T517 ? mem_reg_pc : wb_reg_pc;
  assign T629 = wb_valid;
  assign T630 = T631;
  assign T631 = csr_io_time[6'h20:1'h0];
  assign T632 = io_host_id;
  assign T634 = T68 ? 1'h0 : T635;
  assign T635 = T636 ^ 1'h1;
  assign T636 = wb_reg_valid & wb_ctrl_wxd;
  assign T637 = killm_common & R638;
  assign T639 = div_io_req_ready & T690;
  assign T640 = T103 ? id_ctrl_alu_dw : ex_ctrl_alu_dw;
  assign id_ctrl_alu_dw = T641;
  assign T641 = T644 | T642;
  assign T642 = T643 == 32'h0;
  assign T643 = io_imem_resp_bits_data_0 & 32'h8;
  assign T644 = T645 == 32'h0;
  assign T645 = io_imem_resp_bits_data_0 & 32'h10;
  assign T646 = T103 ? id_ctrl_alu_fn : ex_ctrl_alu_fn;
  assign id_ctrl_alu_fn = T647;
  assign T647 = {T683, T648};
  assign T648 = {T672, T649};
  assign T649 = {T658, T650};
  assign T650 = T653 | T651;
  assign T651 = T652 == 32'h7000;
  assign T652 = io_imem_resp_bits_data_0 & 32'h7044;
  assign T653 = T656 | T654;
  assign T654 = T655 == 32'h1040;
  assign T655 = io_imem_resp_bits_data_0 & 32'h1058;
  assign T656 = T657 == 32'h1010;
  assign T657 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T658 = T661 | T659;
  assign T659 = T660 == 32'h40001010;
  assign T660 = io_imem_resp_bits_data_0 & 32'h40001054;
  assign T661 = T664 | T662;
  assign T662 = T663 == 32'h40000030;
  assign T663 = io_imem_resp_bits_data_0 & 32'h40003034;
  assign T664 = T667 | T665;
  assign T665 = T666 == 32'h6010;
  assign T666 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T667 = T670 | T668;
  assign T668 = T669 == 32'h3010;
  assign T669 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T670 = T671 == 32'h2040;
  assign T671 = io_imem_resp_bits_data_0 & 32'h2058;
  assign T672 = T675 | T673;
  assign T673 = T674 == 32'h4040;
  assign T674 = io_imem_resp_bits_data_0 & 32'h4058;
  assign T675 = T678 | T676;
  assign T676 = T677 == 32'h4010;
  assign T677 = io_imem_resp_bits_data_0 & 32'h5054;
  assign T678 = T681 | T679;
  assign T679 = T680 == 32'h4010;
  assign T680 = io_imem_resp_bits_data_0 & 32'h40004054;
  assign T681 = T682 == 32'h2010;
  assign T682 = io_imem_resp_bits_data_0 & 32'h2054;
  assign T683 = T686 | T684;
  assign T684 = T685 == 32'h40001010;
  assign T685 = io_imem_resp_bits_data_0 & 32'h40003054;
  assign T686 = T687 | T662;
  assign T687 = T212 | T688;
  assign T688 = T689 == 32'h2010;
  assign T689 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T690 = ex_reg_valid & ex_ctrl_div;
  assign T691 = ex_op1;
  assign ex_op1 = T706 ? T705 : T927;
  assign T927 = {T928, T692};
  assign T692 = T694 ? T693 : 40'h0;
  assign T693 = ex_reg_pc;
  assign T694 = ex_ctrl_sel_alu1 == 2'h2;
  assign T695 = T103 ? id_ctrl_sel_alu1 : ex_ctrl_sel_alu1;
  assign id_ctrl_sel_alu1 = T696;
  assign T696 = {T702, T697};
  assign T697 = T698 | T156;
  assign T698 = T699 | T159;
  assign T699 = T161 | T700;
  assign T700 = T701 == 32'h0;
  assign T701 = io_imem_resp_bits_data_0 & 32'h50;
  assign T702 = T703 | T96;
  assign T703 = T704 == 32'h4;
  assign T704 = io_imem_resp_bits_data_0 & 32'h24;
  assign T928 = T929 ? 24'hffffff : 24'h0;
  assign T929 = T692[6'h27:6'h27];
  assign T705 = ex_rs_0;
  assign T706 = ex_ctrl_sel_alu1 == 2'h1;
  assign T707 = ex_op2;
  assign ex_op2 = T806 ? T805 : T930;
  assign T930 = {T936, T708};
  assign T708 = T804 ? ex_imm : T931;
  assign T931 = {T932, T709};
  assign T709 = T710 ? 4'h4 : 4'h0;
  assign T710 = ex_ctrl_sel_alu2 == 2'h1;
  assign T711 = T103 ? id_ctrl_sel_alu2 : ex_ctrl_sel_alu2;
  assign id_ctrl_sel_alu2 = T712;
  assign T712 = {T723, T713};
  assign T713 = T716 | T714;
  assign T714 = T715 == 32'h4050;
  assign T715 = io_imem_resp_bits_data_0 & 32'h4050;
  assign T716 = T717 | T96;
  assign T717 = T718 | T101;
  assign T718 = T721 | T719;
  assign T719 = T720 == 32'h0;
  assign T720 = io_imem_resp_bits_data_0 & 32'h20;
  assign T721 = T722 == 32'h0;
  assign T722 = io_imem_resp_bits_data_0 & 32'h58;
  assign T723 = T726 | T724;
  assign T724 = T725 == 32'h4000;
  assign T725 = io_imem_resp_bits_data_0 & 32'h4008;
  assign T726 = T727 | T156;
  assign T727 = T728 | T159;
  assign T728 = T729 == 32'h0;
  assign T729 = io_imem_resp_bits_data_0 & 32'h48;
  assign T932 = T933 ? 28'hfffffff : 28'h0;
  assign T933 = T709[2'h3:2'h3];
  assign ex_imm = T730;
  assign T730 = {T792, T731};
  assign T731 = {T770, T732};
  assign T732 = {T759, T733};
  assign T733 = T758 ? T757 : T734;
  assign T734 = T756 ? T755 : T735;
  assign T735 = T737 ? T736 : 1'h0;
  assign T736 = ex_reg_inst[4'hf:4'hf];
  assign T737 = ex_ctrl_sel_imm == 3'h5;
  assign T738 = T103 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign id_ctrl_sel_imm = T739;
  assign T739 = {T749, T740};
  assign T740 = {T746, T741};
  assign T741 = T744 | T742;
  assign T742 = T743 == 32'h40;
  assign T743 = io_imem_resp_bits_data_0 & 32'h44;
  assign T744 = T745 == 32'h8;
  assign T745 = io_imem_resp_bits_data_0 & 32'h18;
  assign T746 = T747 | T744;
  assign T747 = T748 == 32'h4;
  assign T748 = io_imem_resp_bits_data_0 & 32'h44;
  assign T749 = T752 | T750;
  assign T750 = T751 == 32'h10;
  assign T751 = io_imem_resp_bits_data_0 & 32'h14;
  assign T752 = T753 | T238;
  assign T753 = T754 == 32'h0;
  assign T754 = io_imem_resp_bits_data_0 & 32'h24;
  assign T755 = ex_reg_inst[5'h14:5'h14];
  assign T756 = ex_ctrl_sel_imm == 3'h4;
  assign T757 = ex_reg_inst[3'h7:3'h7];
  assign T758 = ex_ctrl_sel_imm == 3'h0;
  assign T759 = T769 ? 4'h0 : T760;
  assign T760 = T766 ? T765 : T761;
  assign T761 = T764 ? T763 : T762;
  assign T762 = ex_reg_inst[5'h18:5'h15];
  assign T763 = ex_reg_inst[5'h13:5'h10];
  assign T764 = ex_ctrl_sel_imm == 3'h5;
  assign T765 = ex_reg_inst[4'hb:4'h8];
  assign T766 = T768 | T767;
  assign T767 = ex_ctrl_sel_imm == 3'h1;
  assign T768 = ex_ctrl_sel_imm == 3'h0;
  assign T769 = ex_ctrl_sel_imm == 3'h2;
  assign T770 = {T776, T771};
  assign T771 = T773 ? 6'h0 : T772;
  assign T772 = ex_reg_inst[5'h1e:5'h19];
  assign T773 = T775 | T774;
  assign T774 = ex_ctrl_sel_imm == 3'h5;
  assign T775 = ex_ctrl_sel_imm == 3'h2;
  assign T776 = T789 ? 1'h0 : T777;
  assign T777 = T788 ? T786 : T778;
  assign T778 = T785 ? T783 : T779;
  assign T779 = T782 ? 1'h0 : T780;
  assign T780 = T781;
  assign T781 = ex_reg_inst[5'h1f:5'h1f];
  assign T782 = ex_ctrl_sel_imm == 3'h5;
  assign T783 = T784;
  assign T784 = ex_reg_inst[3'h7:3'h7];
  assign T785 = ex_ctrl_sel_imm == 3'h1;
  assign T786 = T787;
  assign T787 = ex_reg_inst[5'h14:5'h14];
  assign T788 = ex_ctrl_sel_imm == 3'h3;
  assign T789 = T791 | T790;
  assign T790 = ex_ctrl_sel_imm == 3'h5;
  assign T791 = ex_ctrl_sel_imm == 3'h2;
  assign T792 = {T779, T793};
  assign T793 = {T800, T794};
  assign T794 = T797 ? T934 : T795;
  assign T795 = T796;
  assign T796 = ex_reg_inst[5'h13:4'hc];
  assign T934 = T779 ? 8'hff : 8'h0;
  assign T797 = T799 & T798;
  assign T798 = ex_ctrl_sel_imm != 3'h3;
  assign T799 = ex_ctrl_sel_imm != 3'h2;
  assign T800 = T803 ? T801 : T935;
  assign T935 = T779 ? 11'h7ff : 11'h0;
  assign T801 = T802;
  assign T802 = ex_reg_inst[5'h1e:5'h14];
  assign T803 = ex_ctrl_sel_imm == 3'h2;
  assign T804 = ex_ctrl_sel_alu2 == 2'h3;
  assign T936 = T937 ? 32'hffffffff : 32'h0;
  assign T937 = T708[5'h1f:5'h1f];
  assign T805 = ex_rs_1;
  assign T806 = ex_ctrl_sel_alu2 == 2'h2;
  assign T807 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T271 ? mem_reg_cause : T938;
  assign T938 = {61'h0, T808};
  assign T808 = T270 ? 3'h0 : T809;
  assign T809 = T267 ? 3'h6 : T810;
  assign T810 = T264 ? 3'h4 : T811;
  assign T811 = T261 ? 3'h7 : 3'h5;
  assign T812 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T275 ? ex_reg_cause : 64'h2;
  assign T813 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : T939;
  assign T939 = {62'h0, T814};
  assign T814 = io_imem_resp_bits_xcpt_if ? 2'h1 : 2'h2;
  assign T815 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign T816 = wb_reg_inst[5'h1f:5'h14];
  assign io_rocc_exception = T817;
  assign T817 = wb_xcpt & T818;
  assign T818 = csr_io_status_xs != 2'h0;
  assign io_rocc_s = T819;
  assign T819 = csr_io_status_prv != 2'h0;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T820 = T826 ? mem_reg_rs2 : wb_reg_rs2;
  assign T821 = T822 ? ex_rs_1 : mem_reg_rs2;
  assign T822 = T516 & T823;
  assign T823 = ex_ctrl_rxs2 & T824;
  assign T824 = ex_ctrl_mem | ex_ctrl_rocc;
  assign T825 = T103 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign T826 = T517 & mem_ctrl_rocc;
  assign io_rocc_cmd_bits_rs1 = bypass_mux_2;
  assign io_rocc_cmd_bits_inst_opcode = T827;
  assign T827 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T828;
  assign T828 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T829;
  assign T829 = wb_reg_inst[4'hc:4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T830;
  assign T830 = wb_reg_inst[4'hd:4'hd];
  assign io_rocc_cmd_bits_inst_xd = T831;
  assign T831 = wb_reg_inst[4'he:4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T832;
  assign T832 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T833;
  assign T833 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T834;
  assign T834 = wb_reg_inst[5'h1f:5'h19];
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign wb_rocc_val = T836 & T835;
  assign T835 = replay_wb_common ^ 1'h1;
  assign T836 = wb_reg_valid & wb_ctrl_rocc;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = T837;
  assign T837 = T838 & id_ctrl_fp;
  assign T838 = ctrl_killd ^ 1'h1;
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass;
  assign io_fpu_dmem_resp_tag = dmem_resp_waddr;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_val = T839;
  assign T839 = dmem_resp_valid & dmem_resp_fpu;
  assign dmem_resp_fpu = T840;
  assign T840 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data_0;
  assign io_ptw_status_ie = csr_io_status_ie;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_ie1 = csr_io_status_ie1;
  assign io_ptw_status_prv1 = csr_io_status_prv1;
  assign io_ptw_status_ie2 = csr_io_status_ie2;
  assign io_ptw_status_prv2 = csr_io_status_prv2;
  assign io_ptw_status_ie3 = csr_io_status_ie3;
  assign io_ptw_status_prv3 = csr_io_status_prv3;
  assign io_ptw_status_fs = csr_io_status_fs;
  assign io_ptw_status_xs = csr_io_status_xs;
  assign io_ptw_status_mprv = csr_io_status_mprv;
  assign io_ptw_status_vm = csr_io_status_vm;
  assign io_ptw_status_zero1 = csr_io_status_zero1;
  assign io_ptw_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_ptw_status_zero2 = csr_io_status_zero2;
  assign io_ptw_status_sd = csr_io_status_sd;
  assign io_ptw_invalidate = csr_io_fatc;
  assign io_ptw_ptbr = csr_io_ptbr;
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_dmem_req_bits_data = T841;
  assign T841 = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_kill = T842;
  assign T842 = killm_common | mem_xcpt;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_tag = T940;
  assign T940 = {3'h0, T843};
  assign T843 = {ex_waddr, ex_ctrl_fp};
  assign io_dmem_req_bits_addr = T844;
  assign T844 = T845;
  assign T845 = {T847, T846};
  assign T846 = alu_io_adder_out[6'h26:1'h0];
  assign T847 = T860 ? T859 : T848;
  assign T848 = T853 ? T851 : T849;
  assign T849 = T850[1'h0:1'h0];
  assign T850 = alu_io_adder_out[6'h27:6'h26];
  assign T851 = T852 == 2'h3;
  assign T852 = T850;
  assign T853 = T857 | T854;
  assign T854 = T855 == 26'h3fffffe;
  assign T855 = T856;
  assign T856 = ex_rs_0 >> 6'h26;
  assign T857 = T858 == 26'h3ffffff;
  assign T858 = T856;
  assign T859 = T850 != 2'h0;
  assign T860 = T862 | T861;
  assign T861 = T856 == 26'h1;
  assign T862 = T856 == 26'h0;
  assign io_dmem_req_valid = T863;
  assign T863 = ex_reg_valid & ex_ctrl_mem;
  assign io_imem_invalidate = T864;
  assign T864 = wb_reg_valid & wb_ctrl_fence_i;
  assign T865 = T517 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign T866 = T516 ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign T867 = T103 ? id_ctrl_fence_i : ex_ctrl_fence_i;
  assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_returnAddr = T941;
  assign T941 = mem_int_wdata[6'h26:1'h0];
  assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
  assign io_imem_ras_update_bits_isCall = T868;
  assign T868 = mem_ctrl_wxd & T869;
  assign T869 = mem_waddr[1'h0:1'h0];
  assign io_imem_ras_update_valid = T870;
  assign T870 = T872 & T871;
  assign T871 = take_pc_wb ^ 1'h1;
  assign T872 = T874 & T873;
  assign T873 = mem_npc_misaligned ^ 1'h1;
  assign T874 = mem_reg_valid & io_imem_btb_update_bits_isJump;
  assign io_imem_bht_update_bits_mispredict = mem_wrong_npc;
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_pc = T942;
  assign T942 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_bht_update_valid = T875;
  assign T875 = T877 & T876;
  assign T876 = take_pc_wb ^ 1'h1;
  assign T877 = mem_reg_valid & mem_ctrl_branch;
  assign io_imem_btb_update_bits_br_pc = T943;
  assign T943 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_isReturn = T878;
  assign T878 = mem_ctrl_jalr & T879;
  assign T879 = 5'h1 == T880;
  assign T880 = T881 & 5'h19;
  assign T881 = mem_reg_inst[5'h13:4'hf];
  assign io_imem_btb_update_bits_isJump = T882;
  assign T882 = mem_ctrl_jal | mem_ctrl_jalr;
  assign io_imem_btb_update_bits_target = T944;
  assign T944 = io_imem_req_bits_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_pc = T945;
  assign T945 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T883 = T886 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T884 = T885 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T885 = T103 & io_imem_btb_resp_valid;
  assign T886 = T516 & ex_reg_btb_hit;
  assign T887 = T103 ? io_imem_btb_resp_valid : ex_reg_btb_hit;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign T888 = T886 ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign T889 = T885 ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T890 = T886 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T891 = T885 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T892 = T886 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T893 = T885 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign T894 = T886 ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign T895 = T885 ? io_imem_btb_resp_bits_bridx : ex_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign T896 = T886 ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign T897 = T885 ? io_imem_btb_resp_bits_mask : ex_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T898 = T886 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T899 = T885 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T900 = T516 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T901;
  assign T901 = T903 & T902;
  assign T902 = take_pc_wb ^ 1'h1;
  assign T903 = T907 & T904;
  assign T904 = T905 | mem_ctrl_jal;
  assign T905 = T906 | mem_ctrl_jalr;
  assign T906 = mem_ctrl_branch & mem_br_taken;
  assign T907 = T908 & mem_wrong_npc;
  assign T908 = mem_reg_valid & T909;
  assign T909 = mem_npc_misaligned ^ 1'h1;
  assign io_imem_resp_ready = T910;
  assign T910 = T911 | csr_io_interrupt;
  assign T911 = ctrl_stalld ^ 1'h1;
  assign io_imem_req_bits_pc = T912;
  assign T912 = T913;
  assign T913 = T915 ? csr_io_evec : T914;
  assign T914 = replay_wb ? wb_reg_pc : mem_npc;
  assign T915 = wb_xcpt | csr_io_eret;
  assign io_imem_req_valid = take_pc;
  assign io_host_debug_stats_csr = csr_io_host_debug_stats_csr;
  assign io_host_ipi_rep_ready = csr_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = csr_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = csr_io_host_ipi_req_valid;
  assign io_host_csr_resp_bits = csr_io_host_csr_resp_bits;
  assign io_host_csr_resp_valid = csr_io_host_csr_resp_valid;
  assign io_host_csr_req_ready = csr_io_host_csr_req_ready;
  CSRFile csr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_csr_req_ready( csr_io_host_csr_req_ready ),
       .io_host_csr_req_valid( io_host_csr_req_valid ),
       .io_host_csr_req_bits_rw( io_host_csr_req_bits_rw ),
       .io_host_csr_req_bits_addr( io_host_csr_req_bits_addr ),
       .io_host_csr_req_bits_data( io_host_csr_req_bits_data ),
       .io_host_csr_resp_ready( io_host_csr_resp_ready ),
       .io_host_csr_resp_valid( csr_io_host_csr_resp_valid ),
       .io_host_csr_resp_bits( csr_io_host_csr_resp_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( csr_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( csr_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( csr_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_csr( csr_io_host_debug_stats_csr ),
       .io_rw_addr( T816 ),
       .io_rw_cmd( T815 ),
       .io_rw_rdata( csr_io_rw_rdata ),
       .io_rw_wdata( bypass_mux_2 ),
       .io_csr_replay( csr_io_csr_replay ),
       .io_csr_stall( csr_io_csr_stall ),
       .io_csr_xcpt( csr_io_csr_xcpt ),
       .io_eret( csr_io_eret ),
       .io_status_sd( csr_io_status_sd ),
       .io_status_zero2( csr_io_status_zero2 ),
       .io_status_sd_rv32( csr_io_status_sd_rv32 ),
       .io_status_zero1( csr_io_status_zero1 ),
       .io_status_vm( csr_io_status_vm ),
       .io_status_mprv( csr_io_status_mprv ),
       .io_status_xs( csr_io_status_xs ),
       .io_status_fs( csr_io_status_fs ),
       .io_status_prv3( csr_io_status_prv3 ),
       .io_status_ie3( csr_io_status_ie3 ),
       .io_status_prv2( csr_io_status_prv2 ),
       .io_status_ie2( csr_io_status_ie2 ),
       .io_status_prv1( csr_io_status_prv1 ),
       .io_status_ie1( csr_io_status_ie1 ),
       .io_status_prv( csr_io_status_prv ),
       .io_status_ie( csr_io_status_ie ),
       .io_ptbr( csr_io_ptbr ),
       .io_evec( csr_io_evec ),
       .io_exception( wb_reg_xcpt ),
       .io_retire( wb_valid ),
       .io_uarch_counters_15( 1'h0 ),
       .io_uarch_counters_14( 1'h0 ),
       .io_uarch_counters_13( 1'h0 ),
       .io_uarch_counters_12( 1'h0 ),
       .io_uarch_counters_11( 1'h0 ),
       .io_uarch_counters_10( 1'h0 ),
       .io_uarch_counters_9( 1'h0 ),
       .io_uarch_counters_8( 1'h0 ),
       .io_uarch_counters_7( 1'h0 ),
       .io_uarch_counters_6( 1'h0 ),
       .io_uarch_counters_5( 1'h0 ),
       .io_uarch_counters_4( 1'h0 ),
       .io_uarch_counters_3( 1'h0 ),
       .io_uarch_counters_2( 1'h0 ),
       .io_uarch_counters_1( 1'h0 ),
       .io_uarch_counters_0( 1'h0 ),
       .io_cause( wb_reg_cause ),
       .io_pc( wb_reg_pc ),
       .io_fatc( csr_io_fatc ),
       .io_time( csr_io_time ),
       .io_fcsr_rm( csr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_word_bypass(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_invalidate_lr( io_rocc_mem_invalidate_lr ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_addr_block( io_rocc_imem_acquire_bits_addr_block ),
       .io_rocc_imem_acquire_bits_client_xact_id( io_rocc_imem_acquire_bits_client_xact_id ),
       .io_rocc_imem_acquire_bits_addr_beat( io_rocc_imem_acquire_bits_addr_beat ),
       .io_rocc_imem_acquire_bits_is_builtin_type( io_rocc_imem_acquire_bits_is_builtin_type ),
       .io_rocc_imem_acquire_bits_a_type( io_rocc_imem_acquire_bits_a_type ),
       .io_rocc_imem_acquire_bits_union( io_rocc_imem_acquire_bits_union ),
       .io_rocc_imem_acquire_bits_data( io_rocc_imem_acquire_bits_data ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_addr_beat(  )
       //.io_rocc_imem_grant_bits_client_xact_id(  )
       //.io_rocc_imem_grant_bits_manager_xact_id(  )
       //.io_rocc_imem_grant_bits_is_builtin_type(  )
       //.io_rocc_imem_grant_bits_g_type(  )
       //.io_rocc_imem_grant_bits_data(  )
       //.io_rocc_dmem_0_acquire_ready(  )
       .io_rocc_dmem_0_acquire_valid( io_rocc_dmem_0_acquire_valid ),
       .io_rocc_dmem_0_acquire_bits_addr_block( io_rocc_dmem_0_acquire_bits_addr_block ),
       .io_rocc_dmem_0_acquire_bits_client_xact_id( io_rocc_dmem_0_acquire_bits_client_xact_id ),
       .io_rocc_dmem_0_acquire_bits_addr_beat( io_rocc_dmem_0_acquire_bits_addr_beat ),
       .io_rocc_dmem_0_acquire_bits_is_builtin_type( io_rocc_dmem_0_acquire_bits_is_builtin_type ),
       .io_rocc_dmem_0_acquire_bits_a_type( io_rocc_dmem_0_acquire_bits_a_type ),
       .io_rocc_dmem_0_acquire_bits_union( io_rocc_dmem_0_acquire_bits_union ),
       .io_rocc_dmem_0_acquire_bits_data( io_rocc_dmem_0_acquire_bits_data ),
       .io_rocc_dmem_0_grant_ready( io_rocc_dmem_0_grant_ready ),
       //.io_rocc_dmem_0_grant_valid(  )
       //.io_rocc_dmem_0_grant_bits_addr_beat(  )
       //.io_rocc_dmem_0_grant_bits_client_xact_id(  )
       //.io_rocc_dmem_0_grant_bits_manager_xact_id(  )
       //.io_rocc_dmem_0_grant_bits_is_builtin_type(  )
       //.io_rocc_dmem_0_grant_bits_g_type(  )
       //.io_rocc_dmem_0_grant_bits_data(  )
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits_addr( io_rocc_iptw_req_bits_addr ),
       .io_rocc_iptw_req_bits_prv( io_rocc_iptw_req_bits_prv ),
       .io_rocc_iptw_req_bits_store( io_rocc_iptw_req_bits_store ),
       .io_rocc_iptw_req_bits_fetch( io_rocc_iptw_req_bits_fetch ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_pte_ppn(  )
       //.io_rocc_iptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_iptw_resp_bits_pte_d(  )
       //.io_rocc_iptw_resp_bits_pte_r(  )
       //.io_rocc_iptw_resp_bits_pte_typ(  )
       //.io_rocc_iptw_resp_bits_pte_v(  )
       //.io_rocc_iptw_status_sd(  )
       //.io_rocc_iptw_status_zero2(  )
       //.io_rocc_iptw_status_sd_rv32(  )
       //.io_rocc_iptw_status_zero1(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_mprv(  )
       //.io_rocc_iptw_status_xs(  )
       //.io_rocc_iptw_status_fs(  )
       //.io_rocc_iptw_status_prv3(  )
       //.io_rocc_iptw_status_ie3(  )
       //.io_rocc_iptw_status_prv2(  )
       //.io_rocc_iptw_status_ie2(  )
       //.io_rocc_iptw_status_prv1(  )
       //.io_rocc_iptw_status_ie1(  )
       //.io_rocc_iptw_status_prv(  )
       //.io_rocc_iptw_status_ie(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits_addr( io_rocc_dptw_req_bits_addr ),
       .io_rocc_dptw_req_bits_prv( io_rocc_dptw_req_bits_prv ),
       .io_rocc_dptw_req_bits_store( io_rocc_dptw_req_bits_store ),
       .io_rocc_dptw_req_bits_fetch( io_rocc_dptw_req_bits_fetch ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_pte_ppn(  )
       //.io_rocc_dptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_dptw_resp_bits_pte_d(  )
       //.io_rocc_dptw_resp_bits_pte_r(  )
       //.io_rocc_dptw_resp_bits_pte_typ(  )
       //.io_rocc_dptw_resp_bits_pte_v(  )
       //.io_rocc_dptw_status_sd(  )
       //.io_rocc_dptw_status_zero2(  )
       //.io_rocc_dptw_status_sd_rv32(  )
       //.io_rocc_dptw_status_zero1(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_mprv(  )
       //.io_rocc_dptw_status_xs(  )
       //.io_rocc_dptw_status_fs(  )
       //.io_rocc_dptw_status_prv3(  )
       //.io_rocc_dptw_status_ie3(  )
       //.io_rocc_dptw_status_prv2(  )
       //.io_rocc_dptw_status_ie2(  )
       //.io_rocc_dptw_status_prv1(  )
       //.io_rocc_dptw_status_ie1(  )
       //.io_rocc_dptw_status_prv(  )
       //.io_rocc_dptw_status_ie(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits_addr( io_rocc_pptw_req_bits_addr ),
       .io_rocc_pptw_req_bits_prv( io_rocc_pptw_req_bits_prv ),
       .io_rocc_pptw_req_bits_store( io_rocc_pptw_req_bits_store ),
       .io_rocc_pptw_req_bits_fetch( io_rocc_pptw_req_bits_fetch ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_pte_ppn(  )
       //.io_rocc_pptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_pptw_resp_bits_pte_d(  )
       //.io_rocc_pptw_resp_bits_pte_r(  )
       //.io_rocc_pptw_resp_bits_pte_typ(  )
       //.io_rocc_pptw_resp_bits_pte_v(  )
       //.io_rocc_pptw_status_sd(  )
       //.io_rocc_pptw_status_zero2(  )
       //.io_rocc_pptw_status_sd_rv32(  )
       //.io_rocc_pptw_status_zero1(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_mprv(  )
       //.io_rocc_pptw_status_xs(  )
       //.io_rocc_pptw_status_fs(  )
       //.io_rocc_pptw_status_prv3(  )
       //.io_rocc_pptw_status_ie3(  )
       //.io_rocc_pptw_status_prv2(  )
       //.io_rocc_pptw_status_ie2(  )
       //.io_rocc_pptw_status_prv1(  )
       //.io_rocc_pptw_status_ie1(  )
       //.io_rocc_pptw_status_prv(  )
       //.io_rocc_pptw_status_ie(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_exception(  )
       .io_interrupt( csr_io_interrupt ),
       .io_interrupt_cause( csr_io_interrupt_cause )
  );
  ALU alu(
       .io_dw( ex_ctrl_alu_dw ),
       .io_fn( ex_ctrl_alu_fn ),
       .io_in2( T707 ),
       .io_in1( T691 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( T690 ),
       .io_req_bits_fn( ex_ctrl_alu_fn ),
       .io_req_bits_dw( ex_ctrl_alu_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( ex_waddr ),
       .io_kill( T637 ),
       .io_resp_ready( T634 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );

  always @(posedge clk) begin
    if(T517) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T516) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data_0;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T39;
    end
    if(reset) begin
      R73 <= 32'h0;
    end else if(T379) begin
      R73 <= T76;
    end else if(ll_wen) begin
      R73 <= T62;
    end
    if(T517) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if(T516) begin
      mem_ctrl_wxd <= ex_ctrl_wxd;
    end
    if(T103) begin
      ex_ctrl_wxd <= id_ctrl_wxd;
    end
    if(T517) begin
      wb_ctrl_rocc <= mem_ctrl_rocc;
    end
    if(T516) begin
      mem_ctrl_rocc <= ex_ctrl_rocc;
    end
    if(T103) begin
      ex_ctrl_rocc <= id_ctrl_rocc;
    end
    wb_reg_replay <= T114;
    wb_reg_xcpt <= T118;
    if(T516) begin
      mem_ctrl_mem <= ex_ctrl_mem;
    end
    if(T103) begin
      ex_ctrl_mem <= id_ctrl_mem;
    end
    mem_reg_valid <= T124;
    ex_reg_valid <= T126;
    if(T103) begin
      ex_reg_load_use <= id_load_use;
    end
    if(T517) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if(T103) begin
      ex_ctrl_div <= id_ctrl_div;
    end
    if(T516) begin
      mem_ctrl_jal <= ex_ctrl_jal;
    end
    if(T103) begin
      ex_ctrl_jal <= id_ctrl_jal;
    end
    if(T516) begin
      bypass_mux_1 <= alu_io_out;
    end
    if(T516) begin
      mem_ctrl_branch <= ex_ctrl_branch;
    end
    if(T103) begin
      ex_ctrl_branch <= id_ctrl_branch;
    end
    if(T516) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T516) begin
      mem_ctrl_jalr <= ex_ctrl_jalr;
    end
    if(T103) begin
      ex_ctrl_jalr <= id_ctrl_jalr;
    end
    if(T516) begin
      mem_reg_flush_pipe <= ex_reg_flush_pipe;
    end
    if(T103) begin
      ex_reg_flush_pipe <= T243;
    end
    mem_reg_xcpt <= T272;
    if(T103) begin
      ex_ctrl_fp <= id_ctrl_fp;
    end
    ex_reg_xcpt <= T276;
    ex_reg_xcpt_interrupt <= T359;
    mem_reg_xcpt_interrupt <= T363;
    if(T516) begin
      mem_ctrl_fp <= ex_ctrl_fp;
    end
    mem_reg_replay <= T368;
    wb_reg_valid <= T371;
    if(T517) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if(T516) begin
      mem_ctrl_div <= ex_ctrl_div;
    end
    if(T517) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if(T516) begin
      mem_ctrl_wfd <= ex_ctrl_wfd;
    end
    if(T103) begin
      ex_ctrl_wfd <= id_ctrl_wfd;
    end
    if(T516) begin
      mem_mem_cmd_bh <= ex_slow_bypass;
    end
    if(T103) begin
      ex_ctrl_mem_type <= id_ctrl_mem_type;
    end
    if(T103) begin
      ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
    end
    if(T516) begin
      mem_ctrl_csr <= ex_ctrl_csr;
    end
    if(T103) begin
      ex_ctrl_csr <= id_csr;
    end else if(T103) begin
      ex_ctrl_csr <= id_ctrl_csr;
    end
    R521 <= R522;
    if(ex_reg_rs_bypass_1) begin
      R522 <= T573;
    end else begin
      R522 <= T523;
    end
    if(T562) begin
      ex_reg_rs_lsb_1 <= T538;
    end else if(T103) begin
      ex_reg_rs_lsb_1 <= T526;
    end
    if (T543)
      T541[T548] <= rf_wdata;
    if(T517) begin
      bypass_mux_2 <= T553;
    end
    if(T517) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if(T562) begin
      ex_reg_rs_msb_1 <= T572;
    end
    if(T103) begin
      ex_reg_rs_bypass_1 <= T565;
    end
    R584 <= R585;
    if(ex_reg_rs_bypass_0) begin
      R585 <= T613;
    end else begin
      R585 <= T586;
    end
    if(T603) begin
      ex_reg_rs_lsb_0 <= T597;
    end else if(T103) begin
      ex_reg_rs_lsb_0 <= T589;
    end
    if(T603) begin
      ex_reg_rs_msb_0 <= T612;
    end
    if(T103) begin
      ex_reg_rs_bypass_0 <= T606;
    end
    if(T517) begin
      wb_reg_pc <= mem_reg_pc;
    end
    R638 <= T639;
    if(T103) begin
      ex_ctrl_alu_dw <= id_ctrl_alu_dw;
    end
    if(T103) begin
      ex_ctrl_alu_fn <= id_ctrl_alu_fn;
    end
    if(T103) begin
      ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
    end
    if(T103) begin
      ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
    end
    if(T103) begin
      ex_ctrl_sel_imm <= id_ctrl_sel_imm;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(T826) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(T822) begin
      mem_reg_rs2 <= ex_rs_1;
    end
    if(T103) begin
      ex_ctrl_rxs2 <= id_ctrl_rxs2;
    end
    if(T517) begin
      wb_ctrl_fence_i <= mem_ctrl_fence_i;
    end
    if(T516) begin
      mem_ctrl_fence_i <= ex_ctrl_fence_i;
    end
    if(T103) begin
      ex_ctrl_fence_i <= id_ctrl_fence_i;
    end
    if(T886) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T885) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(T103) begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T886) begin
      mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
    end
    if(T885) begin
      ex_reg_btb_resp_bht_history <= io_imem_btb_resp_bits_bht_history;
    end
    if(T886) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T885) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T886) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T885) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T886) begin
      mem_reg_btb_resp_bridx <= ex_reg_btb_resp_bridx;
    end
    if(T885) begin
      ex_reg_btb_resp_bridx <= io_imem_btb_resp_bits_bridx;
    end
    if(T886) begin
      mem_reg_btb_resp_mask <= ex_reg_btb_resp_mask;
    end
    if(T885) begin
      ex_reg_btb_resp_mask <= io_imem_btb_resp_bits_mask;
    end
    if(T886) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T885) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T516) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T632, T630, T629, T627, T625, T624, T623, T621, T583, T581, T520, T519, T1);
// synthesis translate_on
`endif
  end
endmodule

module BTB(input clk, input reset,
    input  io_req_valid,
    input [38:0] io_req_bits_addr,
    output io_resp_valid,
    output io_resp_bits_taken,
    output io_resp_bits_mask,
    output io_resp_bits_bridx,
    output[38:0] io_resp_bits_target,
    output[5:0] io_resp_bits_entry,
    output[6:0] io_resp_bits_bht_history,
    output[1:0] io_resp_bits_bht_value,
    input  io_btb_update_valid,
    input  io_btb_update_bits_prediction_valid,
    input  io_btb_update_bits_prediction_bits_taken,
    input  io_btb_update_bits_prediction_bits_mask,
    input  io_btb_update_bits_prediction_bits_bridx,
    input [38:0] io_btb_update_bits_prediction_bits_target,
    input [5:0] io_btb_update_bits_prediction_bits_entry,
    input [6:0] io_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_btb_update_bits_prediction_bits_bht_value,
    input [38:0] io_btb_update_bits_pc,
    input [38:0] io_btb_update_bits_target,
    input  io_btb_update_bits_taken,
    input  io_btb_update_bits_isJump,
    input  io_btb_update_bits_isReturn,
    input [38:0] io_btb_update_bits_br_pc,
    input  io_bht_update_valid,
    input  io_bht_update_bits_prediction_valid,
    input  io_bht_update_bits_prediction_bits_taken,
    input  io_bht_update_bits_prediction_bits_mask,
    input  io_bht_update_bits_prediction_bits_bridx,
    input [38:0] io_bht_update_bits_prediction_bits_target,
    input [5:0] io_bht_update_bits_prediction_bits_entry,
    input [6:0] io_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_bht_update_bits_prediction_bits_bht_value,
    input [38:0] io_bht_update_bits_pc,
    input  io_bht_update_bits_taken,
    input  io_bht_update_bits_mispredict,
    input  io_ras_update_valid,
    input  io_ras_update_bits_isCall,
    input  io_ras_update_bits_isReturn,
    input [38:0] io_ras_update_bits_returnAddr,
    input  io_ras_update_bits_prediction_valid,
    input  io_ras_update_bits_prediction_bits_taken,
    input  io_ras_update_bits_prediction_bits_mask,
    input  io_ras_update_bits_prediction_bits_bridx,
    input [38:0] io_ras_update_bits_prediction_bits_target,
    input [5:0] io_ras_update_bits_prediction_bits_entry,
    input [6:0] io_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_ras_update_bits_prediction_bits_bht_value,
    input  io_invalidate
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg [38:0] R4;
  wire[38:0] T5;
  wire T6;
  reg  R7;
  wire T2288;
  wire[1:0] T8;
  wire[1:0] T9;
  reg [1:0] T10 [127:0];
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[6:0] T22;
  wire[6:0] T23;
  wire[6:0] T24;
  reg [6:0] R25;
  wire[6:0] T26;
  wire[6:0] T27;
  wire[6:0] T28;
  wire[5:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  reg  isJump_61;
  wire T35;
  reg  R36;
  wire T37;
  wire T38;
  wire T39;
  wire[63:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  reg [5:0] nextRepl;
  wire[5:0] T2289;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire T46;
  wire T47;
  wire T48;
  reg [5:0] R49;
  wire[5:0] T50;
  reg  updateHit;
  wire T51;
  wire T52;
  wire[61:0] hits;
  wire[61:0] T53;
  wire[61:0] T54;
  wire[30:0] T55;
  wire[15:0] T56;
  wire[7:0] T57;
  wire[3:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[5:0] T61;
  wire[5:0] pageHit;
  reg [5:0] pageValid;
  wire[5:0] T2290;
  wire[5:0] T62;
  wire[5:0] T63;
  wire[5:0] T64;
  wire[5:0] pageReplEn;
  wire[5:0] tgtPageReplEn;
  wire[5:0] tgtPageRepl;
  wire[5:0] T65;
  wire[5:0] T2291;
  wire T66;
  wire[5:0] T67;
  wire[4:0] T68;
  wire[5:0] idxPageUpdateOH;
  wire[5:0] idxPageRepl;
  wire[5:0] T2292;
  wire[7:0] T69;
  reg [2:0] R70;
  wire[2:0] T2293;
  wire[2:0] T71;
  wire[2:0] T72;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire doPageRepl;
  wire doIdxPageRepl;
  wire[5:0] updatePageHit;
  wire[5:0] T76;
  wire[5:0] T77;
  wire[2:0] T78;
  wire[1:0] T79;
  wire T80;
  wire[26:0] T81;
  reg [38:0] R82;
  wire[38:0] T83;
  wire[26:0] T84;
  reg [26:0] pages [5:0];
  wire[26:0] T85;
  wire[26:0] T86;
  wire[26:0] T87;
  wire[26:0] T88;
  wire T89;
  wire[5:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire[26:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire[26:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[26:0] T103;
  wire[26:0] T104;
  wire[26:0] T105;
  wire[26:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire[26:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire[26:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire[26:0] T120;
  wire T121;
  wire[26:0] T122;
  wire[2:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[26:0] T126;
  wire T127;
  wire[26:0] T128;
  wire T129;
  wire[26:0] T130;
  wire useUpdatePageHit;
  wire samePage;
  wire[26:0] T131;
  wire[26:0] T132;
  wire doTgtPageRepl;
  wire T133;
  wire usePageHit;
  wire[5:0] T134;
  wire[5:0] T135;
  wire T136;
  wire[5:0] idxPageReplEn;
  wire T137;
  wire[5:0] T138;
  wire[5:0] T139;
  wire[2:0] T140;
  wire[1:0] T141;
  wire T142;
  wire[26:0] T143;
  wire[26:0] T144;
  wire T145;
  wire[26:0] T146;
  wire T147;
  wire[26:0] T148;
  wire[2:0] T149;
  wire[1:0] T150;
  wire T151;
  wire[26:0] T152;
  wire T153;
  wire[26:0] T154;
  wire T155;
  wire[26:0] T156;
  wire[5:0] idxPagesOH_0;
  wire[7:0] T157;
  wire[2:0] T158;
  reg [2:0] idxPages [61:0];
  wire[2:0] T159;
  wire[2:0] T2294;
  wire[1:0] T2295;
  wire T2296;
  wire[1:0] T2297;
  wire[1:0] T2298;
  wire[3:0] T2299;
  wire[3:0] T2300;
  wire[1:0] T2301;
  wire[1:0] T2302;
  wire T2303;
  wire T2304;
  wire T160;
  wire T161;
  wire T162;
  wire[5:0] T163;
  wire[5:0] idxPagesOH_1;
  wire[7:0] T164;
  wire[2:0] T165;
  wire[1:0] T166;
  wire T167;
  wire[5:0] T168;
  wire[5:0] idxPagesOH_2;
  wire[7:0] T169;
  wire[2:0] T170;
  wire T171;
  wire[5:0] T172;
  wire[5:0] idxPagesOH_3;
  wire[7:0] T173;
  wire[2:0] T174;
  wire[3:0] T175;
  wire[1:0] T176;
  wire T177;
  wire[5:0] T178;
  wire[5:0] idxPagesOH_4;
  wire[7:0] T179;
  wire[2:0] T180;
  wire T181;
  wire[5:0] T182;
  wire[5:0] idxPagesOH_5;
  wire[7:0] T183;
  wire[2:0] T184;
  wire[1:0] T185;
  wire T186;
  wire[5:0] T187;
  wire[5:0] idxPagesOH_6;
  wire[7:0] T188;
  wire[2:0] T189;
  wire T190;
  wire[5:0] T191;
  wire[5:0] idxPagesOH_7;
  wire[7:0] T192;
  wire[2:0] T193;
  wire[7:0] T194;
  wire[3:0] T195;
  wire[1:0] T196;
  wire T197;
  wire[5:0] T198;
  wire[5:0] idxPagesOH_8;
  wire[7:0] T199;
  wire[2:0] T200;
  wire T201;
  wire[5:0] T202;
  wire[5:0] idxPagesOH_9;
  wire[7:0] T203;
  wire[2:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[5:0] T207;
  wire[5:0] idxPagesOH_10;
  wire[7:0] T208;
  wire[2:0] T209;
  wire T210;
  wire[5:0] T211;
  wire[5:0] idxPagesOH_11;
  wire[7:0] T212;
  wire[2:0] T213;
  wire[3:0] T214;
  wire[1:0] T215;
  wire T216;
  wire[5:0] T217;
  wire[5:0] idxPagesOH_12;
  wire[7:0] T218;
  wire[2:0] T219;
  wire T220;
  wire[5:0] T221;
  wire[5:0] idxPagesOH_13;
  wire[7:0] T222;
  wire[2:0] T223;
  wire[1:0] T224;
  wire T225;
  wire[5:0] T226;
  wire[5:0] idxPagesOH_14;
  wire[7:0] T227;
  wire[2:0] T228;
  wire T229;
  wire[5:0] T230;
  wire[5:0] idxPagesOH_15;
  wire[7:0] T231;
  wire[2:0] T232;
  wire[14:0] T233;
  wire[7:0] T234;
  wire[3:0] T235;
  wire[1:0] T236;
  wire T237;
  wire[5:0] T238;
  wire[5:0] idxPagesOH_16;
  wire[7:0] T239;
  wire[2:0] T240;
  wire T241;
  wire[5:0] T242;
  wire[5:0] idxPagesOH_17;
  wire[7:0] T243;
  wire[2:0] T244;
  wire[1:0] T245;
  wire T246;
  wire[5:0] T247;
  wire[5:0] idxPagesOH_18;
  wire[7:0] T248;
  wire[2:0] T249;
  wire T250;
  wire[5:0] T251;
  wire[5:0] idxPagesOH_19;
  wire[7:0] T252;
  wire[2:0] T253;
  wire[3:0] T254;
  wire[1:0] T255;
  wire T256;
  wire[5:0] T257;
  wire[5:0] idxPagesOH_20;
  wire[7:0] T258;
  wire[2:0] T259;
  wire T260;
  wire[5:0] T261;
  wire[5:0] idxPagesOH_21;
  wire[7:0] T262;
  wire[2:0] T263;
  wire[1:0] T264;
  wire T265;
  wire[5:0] T266;
  wire[5:0] idxPagesOH_22;
  wire[7:0] T267;
  wire[2:0] T268;
  wire T269;
  wire[5:0] T270;
  wire[5:0] idxPagesOH_23;
  wire[7:0] T271;
  wire[2:0] T272;
  wire[6:0] T273;
  wire[3:0] T274;
  wire[1:0] T275;
  wire T276;
  wire[5:0] T277;
  wire[5:0] idxPagesOH_24;
  wire[7:0] T278;
  wire[2:0] T279;
  wire T280;
  wire[5:0] T281;
  wire[5:0] idxPagesOH_25;
  wire[7:0] T282;
  wire[2:0] T283;
  wire[1:0] T284;
  wire T285;
  wire[5:0] T286;
  wire[5:0] idxPagesOH_26;
  wire[7:0] T287;
  wire[2:0] T288;
  wire T289;
  wire[5:0] T290;
  wire[5:0] idxPagesOH_27;
  wire[7:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[1:0] T294;
  wire T295;
  wire[5:0] T296;
  wire[5:0] idxPagesOH_28;
  wire[7:0] T297;
  wire[2:0] T298;
  wire T299;
  wire[5:0] T300;
  wire[5:0] idxPagesOH_29;
  wire[7:0] T301;
  wire[2:0] T302;
  wire T303;
  wire[5:0] T304;
  wire[5:0] idxPagesOH_30;
  wire[7:0] T305;
  wire[2:0] T306;
  wire[30:0] T307;
  wire[15:0] T308;
  wire[7:0] T309;
  wire[3:0] T310;
  wire[1:0] T311;
  wire T312;
  wire[5:0] T313;
  wire[5:0] idxPagesOH_31;
  wire[7:0] T314;
  wire[2:0] T315;
  wire T316;
  wire[5:0] T317;
  wire[5:0] idxPagesOH_32;
  wire[7:0] T318;
  wire[2:0] T319;
  wire[1:0] T320;
  wire T321;
  wire[5:0] T322;
  wire[5:0] idxPagesOH_33;
  wire[7:0] T323;
  wire[2:0] T324;
  wire T325;
  wire[5:0] T326;
  wire[5:0] idxPagesOH_34;
  wire[7:0] T327;
  wire[2:0] T328;
  wire[3:0] T329;
  wire[1:0] T330;
  wire T331;
  wire[5:0] T332;
  wire[5:0] idxPagesOH_35;
  wire[7:0] T333;
  wire[2:0] T334;
  wire T335;
  wire[5:0] T336;
  wire[5:0] idxPagesOH_36;
  wire[7:0] T337;
  wire[2:0] T338;
  wire[1:0] T339;
  wire T340;
  wire[5:0] T341;
  wire[5:0] idxPagesOH_37;
  wire[7:0] T342;
  wire[2:0] T343;
  wire T344;
  wire[5:0] T345;
  wire[5:0] idxPagesOH_38;
  wire[7:0] T346;
  wire[2:0] T347;
  wire[7:0] T348;
  wire[3:0] T349;
  wire[1:0] T350;
  wire T351;
  wire[5:0] T352;
  wire[5:0] idxPagesOH_39;
  wire[7:0] T353;
  wire[2:0] T354;
  wire T355;
  wire[5:0] T356;
  wire[5:0] idxPagesOH_40;
  wire[7:0] T357;
  wire[2:0] T358;
  wire[1:0] T359;
  wire T360;
  wire[5:0] T361;
  wire[5:0] idxPagesOH_41;
  wire[7:0] T362;
  wire[2:0] T363;
  wire T364;
  wire[5:0] T365;
  wire[5:0] idxPagesOH_42;
  wire[7:0] T366;
  wire[2:0] T367;
  wire[3:0] T368;
  wire[1:0] T369;
  wire T370;
  wire[5:0] T371;
  wire[5:0] idxPagesOH_43;
  wire[7:0] T372;
  wire[2:0] T373;
  wire T374;
  wire[5:0] T375;
  wire[5:0] idxPagesOH_44;
  wire[7:0] T376;
  wire[2:0] T377;
  wire[1:0] T378;
  wire T379;
  wire[5:0] T380;
  wire[5:0] idxPagesOH_45;
  wire[7:0] T381;
  wire[2:0] T382;
  wire T383;
  wire[5:0] T384;
  wire[5:0] idxPagesOH_46;
  wire[7:0] T385;
  wire[2:0] T386;
  wire[14:0] T387;
  wire[7:0] T388;
  wire[3:0] T389;
  wire[1:0] T390;
  wire T391;
  wire[5:0] T392;
  wire[5:0] idxPagesOH_47;
  wire[7:0] T393;
  wire[2:0] T394;
  wire T395;
  wire[5:0] T396;
  wire[5:0] idxPagesOH_48;
  wire[7:0] T397;
  wire[2:0] T398;
  wire[1:0] T399;
  wire T400;
  wire[5:0] T401;
  wire[5:0] idxPagesOH_49;
  wire[7:0] T402;
  wire[2:0] T403;
  wire T404;
  wire[5:0] T405;
  wire[5:0] idxPagesOH_50;
  wire[7:0] T406;
  wire[2:0] T407;
  wire[3:0] T408;
  wire[1:0] T409;
  wire T410;
  wire[5:0] T411;
  wire[5:0] idxPagesOH_51;
  wire[7:0] T412;
  wire[2:0] T413;
  wire T414;
  wire[5:0] T415;
  wire[5:0] idxPagesOH_52;
  wire[7:0] T416;
  wire[2:0] T417;
  wire[1:0] T418;
  wire T419;
  wire[5:0] T420;
  wire[5:0] idxPagesOH_53;
  wire[7:0] T421;
  wire[2:0] T422;
  wire T423;
  wire[5:0] T424;
  wire[5:0] idxPagesOH_54;
  wire[7:0] T425;
  wire[2:0] T426;
  wire[6:0] T427;
  wire[3:0] T428;
  wire[1:0] T429;
  wire T430;
  wire[5:0] T431;
  wire[5:0] idxPagesOH_55;
  wire[7:0] T432;
  wire[2:0] T433;
  wire T434;
  wire[5:0] T435;
  wire[5:0] idxPagesOH_56;
  wire[7:0] T436;
  wire[2:0] T437;
  wire[1:0] T438;
  wire T439;
  wire[5:0] T440;
  wire[5:0] idxPagesOH_57;
  wire[7:0] T441;
  wire[2:0] T442;
  wire T443;
  wire[5:0] T444;
  wire[5:0] idxPagesOH_58;
  wire[7:0] T445;
  wire[2:0] T446;
  wire[2:0] T447;
  wire[1:0] T448;
  wire T449;
  wire[5:0] T450;
  wire[5:0] idxPagesOH_59;
  wire[7:0] T451;
  wire[2:0] T452;
  wire T453;
  wire[5:0] T454;
  wire[5:0] idxPagesOH_60;
  wire[7:0] T455;
  wire[2:0] T456;
  wire T457;
  wire[5:0] T458;
  wire[5:0] idxPagesOH_61;
  wire[7:0] T459;
  wire[2:0] T460;
  wire[61:0] T461;
  wire[61:0] T462;
  wire[61:0] T463;
  wire[30:0] T464;
  wire[15:0] T465;
  wire[7:0] T466;
  wire[3:0] T467;
  wire[1:0] T468;
  wire T469;
  wire[11:0] T470;
  wire[11:0] T471;
  reg [11:0] idxs [61:0];
  wire[11:0] T472;
  wire[11:0] T2305;
  wire T473;
  wire T474;
  wire T475;
  wire[11:0] T476;
  wire[1:0] T477;
  wire T478;
  wire[11:0] T479;
  wire T480;
  wire[11:0] T481;
  wire[3:0] T482;
  wire[1:0] T483;
  wire T484;
  wire[11:0] T485;
  wire T486;
  wire[11:0] T487;
  wire[1:0] T488;
  wire T489;
  wire[11:0] T490;
  wire T491;
  wire[11:0] T492;
  wire[7:0] T493;
  wire[3:0] T494;
  wire[1:0] T495;
  wire T496;
  wire[11:0] T497;
  wire T498;
  wire[11:0] T499;
  wire[1:0] T500;
  wire T501;
  wire[11:0] T502;
  wire T503;
  wire[11:0] T504;
  wire[3:0] T505;
  wire[1:0] T506;
  wire T507;
  wire[11:0] T508;
  wire T509;
  wire[11:0] T510;
  wire[1:0] T511;
  wire T512;
  wire[11:0] T513;
  wire T514;
  wire[11:0] T515;
  wire[14:0] T516;
  wire[7:0] T517;
  wire[3:0] T518;
  wire[1:0] T519;
  wire T520;
  wire[11:0] T521;
  wire T522;
  wire[11:0] T523;
  wire[1:0] T524;
  wire T525;
  wire[11:0] T526;
  wire T527;
  wire[11:0] T528;
  wire[3:0] T529;
  wire[1:0] T530;
  wire T531;
  wire[11:0] T532;
  wire T533;
  wire[11:0] T534;
  wire[1:0] T535;
  wire T536;
  wire[11:0] T537;
  wire T538;
  wire[11:0] T539;
  wire[6:0] T540;
  wire[3:0] T541;
  wire[1:0] T542;
  wire T543;
  wire[11:0] T544;
  wire T545;
  wire[11:0] T546;
  wire[1:0] T547;
  wire T548;
  wire[11:0] T549;
  wire T550;
  wire[11:0] T551;
  wire[2:0] T552;
  wire[1:0] T553;
  wire T554;
  wire[11:0] T555;
  wire T556;
  wire[11:0] T557;
  wire T558;
  wire[11:0] T559;
  wire[30:0] T560;
  wire[15:0] T561;
  wire[7:0] T562;
  wire[3:0] T563;
  wire[1:0] T564;
  wire T565;
  wire[11:0] T566;
  wire T567;
  wire[11:0] T568;
  wire[1:0] T569;
  wire T570;
  wire[11:0] T571;
  wire T572;
  wire[11:0] T573;
  wire[3:0] T574;
  wire[1:0] T575;
  wire T576;
  wire[11:0] T577;
  wire T578;
  wire[11:0] T579;
  wire[1:0] T580;
  wire T581;
  wire[11:0] T582;
  wire T583;
  wire[11:0] T584;
  wire[7:0] T585;
  wire[3:0] T586;
  wire[1:0] T587;
  wire T588;
  wire[11:0] T589;
  wire T590;
  wire[11:0] T591;
  wire[1:0] T592;
  wire T593;
  wire[11:0] T594;
  wire T595;
  wire[11:0] T596;
  wire[3:0] T597;
  wire[1:0] T598;
  wire T599;
  wire[11:0] T600;
  wire T601;
  wire[11:0] T602;
  wire[1:0] T603;
  wire T604;
  wire[11:0] T605;
  wire T606;
  wire[11:0] T607;
  wire[14:0] T608;
  wire[7:0] T609;
  wire[3:0] T610;
  wire[1:0] T611;
  wire T612;
  wire[11:0] T613;
  wire T614;
  wire[11:0] T615;
  wire[1:0] T616;
  wire T617;
  wire[11:0] T618;
  wire T619;
  wire[11:0] T620;
  wire[3:0] T621;
  wire[1:0] T622;
  wire T623;
  wire[11:0] T624;
  wire T625;
  wire[11:0] T626;
  wire[1:0] T627;
  wire T628;
  wire[11:0] T629;
  wire T630;
  wire[11:0] T631;
  wire[6:0] T632;
  wire[3:0] T633;
  wire[1:0] T634;
  wire T635;
  wire[11:0] T636;
  wire T637;
  wire[11:0] T638;
  wire[1:0] T639;
  wire T640;
  wire[11:0] T641;
  wire T642;
  wire[11:0] T643;
  wire[2:0] T644;
  wire[1:0] T645;
  wire T646;
  wire[11:0] T647;
  wire T648;
  wire[11:0] T649;
  wire T650;
  wire[11:0] T651;
  reg [61:0] idxValid;
  wire[61:0] T2306;
  wire[63:0] T2307;
  wire[63:0] T652;
  wire[63:0] T653;
  wire[63:0] T2308;
  wire[63:0] T654;
  wire[63:0] T655;
  wire[63:0] T2309;
  wire[61:0] T656;
  wire[61:0] T657;
  wire[61:0] T658;
  wire[61:0] T659;
  wire[30:0] T660;
  wire[15:0] T661;
  wire[7:0] T662;
  wire[3:0] T663;
  wire[1:0] T664;
  wire T665;
  wire[5:0] T666;
  wire[5:0] T667;
  wire[5:0] tgtPagesOH_0;
  wire[7:0] T668;
  wire[2:0] T669;
  reg [2:0] tgtPages [61:0];
  wire[2:0] T670;
  wire[2:0] T2310;
  wire[1:0] T2311;
  wire T2312;
  wire[1:0] T2313;
  wire[1:0] T2314;
  wire[3:0] T2315;
  wire[3:0] T2316;
  wire[5:0] T671;
  wire[1:0] T2317;
  wire[1:0] T2318;
  wire T2319;
  wire T2320;
  wire T672;
  wire T673;
  wire T674;
  wire[5:0] T675;
  wire[5:0] T676;
  wire[5:0] tgtPagesOH_1;
  wire[7:0] T677;
  wire[2:0] T678;
  wire[1:0] T679;
  wire T680;
  wire[5:0] T681;
  wire[5:0] T682;
  wire[5:0] tgtPagesOH_2;
  wire[7:0] T683;
  wire[2:0] T684;
  wire T685;
  wire[5:0] T686;
  wire[5:0] T687;
  wire[5:0] tgtPagesOH_3;
  wire[7:0] T688;
  wire[2:0] T689;
  wire[3:0] T690;
  wire[1:0] T691;
  wire T692;
  wire[5:0] T693;
  wire[5:0] T694;
  wire[5:0] tgtPagesOH_4;
  wire[7:0] T695;
  wire[2:0] T696;
  wire T697;
  wire[5:0] T698;
  wire[5:0] T699;
  wire[5:0] tgtPagesOH_5;
  wire[7:0] T700;
  wire[2:0] T701;
  wire[1:0] T702;
  wire T703;
  wire[5:0] T704;
  wire[5:0] T705;
  wire[5:0] tgtPagesOH_6;
  wire[7:0] T706;
  wire[2:0] T707;
  wire T708;
  wire[5:0] T709;
  wire[5:0] T710;
  wire[5:0] tgtPagesOH_7;
  wire[7:0] T711;
  wire[2:0] T712;
  wire[7:0] T713;
  wire[3:0] T714;
  wire[1:0] T715;
  wire T716;
  wire[5:0] T717;
  wire[5:0] T718;
  wire[5:0] tgtPagesOH_8;
  wire[7:0] T719;
  wire[2:0] T720;
  wire T721;
  wire[5:0] T722;
  wire[5:0] T723;
  wire[5:0] tgtPagesOH_9;
  wire[7:0] T724;
  wire[2:0] T725;
  wire[1:0] T726;
  wire T727;
  wire[5:0] T728;
  wire[5:0] T729;
  wire[5:0] tgtPagesOH_10;
  wire[7:0] T730;
  wire[2:0] T731;
  wire T732;
  wire[5:0] T733;
  wire[5:0] T734;
  wire[5:0] tgtPagesOH_11;
  wire[7:0] T735;
  wire[2:0] T736;
  wire[3:0] T737;
  wire[1:0] T738;
  wire T739;
  wire[5:0] T740;
  wire[5:0] T741;
  wire[5:0] tgtPagesOH_12;
  wire[7:0] T742;
  wire[2:0] T743;
  wire T744;
  wire[5:0] T745;
  wire[5:0] T746;
  wire[5:0] tgtPagesOH_13;
  wire[7:0] T747;
  wire[2:0] T748;
  wire[1:0] T749;
  wire T750;
  wire[5:0] T751;
  wire[5:0] T752;
  wire[5:0] tgtPagesOH_14;
  wire[7:0] T753;
  wire[2:0] T754;
  wire T755;
  wire[5:0] T756;
  wire[5:0] T757;
  wire[5:0] tgtPagesOH_15;
  wire[7:0] T758;
  wire[2:0] T759;
  wire[14:0] T760;
  wire[7:0] T761;
  wire[3:0] T762;
  wire[1:0] T763;
  wire T764;
  wire[5:0] T765;
  wire[5:0] T766;
  wire[5:0] tgtPagesOH_16;
  wire[7:0] T767;
  wire[2:0] T768;
  wire T769;
  wire[5:0] T770;
  wire[5:0] T771;
  wire[5:0] tgtPagesOH_17;
  wire[7:0] T772;
  wire[2:0] T773;
  wire[1:0] T774;
  wire T775;
  wire[5:0] T776;
  wire[5:0] T777;
  wire[5:0] tgtPagesOH_18;
  wire[7:0] T778;
  wire[2:0] T779;
  wire T780;
  wire[5:0] T781;
  wire[5:0] T782;
  wire[5:0] tgtPagesOH_19;
  wire[7:0] T783;
  wire[2:0] T784;
  wire[3:0] T785;
  wire[1:0] T786;
  wire T787;
  wire[5:0] T788;
  wire[5:0] T789;
  wire[5:0] tgtPagesOH_20;
  wire[7:0] T790;
  wire[2:0] T791;
  wire T792;
  wire[5:0] T793;
  wire[5:0] T794;
  wire[5:0] tgtPagesOH_21;
  wire[7:0] T795;
  wire[2:0] T796;
  wire[1:0] T797;
  wire T798;
  wire[5:0] T799;
  wire[5:0] T800;
  wire[5:0] tgtPagesOH_22;
  wire[7:0] T801;
  wire[2:0] T802;
  wire T803;
  wire[5:0] T804;
  wire[5:0] T805;
  wire[5:0] tgtPagesOH_23;
  wire[7:0] T806;
  wire[2:0] T807;
  wire[6:0] T808;
  wire[3:0] T809;
  wire[1:0] T810;
  wire T811;
  wire[5:0] T812;
  wire[5:0] T813;
  wire[5:0] tgtPagesOH_24;
  wire[7:0] T814;
  wire[2:0] T815;
  wire T816;
  wire[5:0] T817;
  wire[5:0] T818;
  wire[5:0] tgtPagesOH_25;
  wire[7:0] T819;
  wire[2:0] T820;
  wire[1:0] T821;
  wire T822;
  wire[5:0] T823;
  wire[5:0] T824;
  wire[5:0] tgtPagesOH_26;
  wire[7:0] T825;
  wire[2:0] T826;
  wire T827;
  wire[5:0] T828;
  wire[5:0] T829;
  wire[5:0] tgtPagesOH_27;
  wire[7:0] T830;
  wire[2:0] T831;
  wire[2:0] T832;
  wire[1:0] T833;
  wire T834;
  wire[5:0] T835;
  wire[5:0] T836;
  wire[5:0] tgtPagesOH_28;
  wire[7:0] T837;
  wire[2:0] T838;
  wire T839;
  wire[5:0] T840;
  wire[5:0] T841;
  wire[5:0] tgtPagesOH_29;
  wire[7:0] T842;
  wire[2:0] T843;
  wire T844;
  wire[5:0] T845;
  wire[5:0] T846;
  wire[5:0] tgtPagesOH_30;
  wire[7:0] T847;
  wire[2:0] T848;
  wire[30:0] T849;
  wire[15:0] T850;
  wire[7:0] T851;
  wire[3:0] T852;
  wire[1:0] T853;
  wire T854;
  wire[5:0] T855;
  wire[5:0] T856;
  wire[5:0] tgtPagesOH_31;
  wire[7:0] T857;
  wire[2:0] T858;
  wire T859;
  wire[5:0] T860;
  wire[5:0] T861;
  wire[5:0] tgtPagesOH_32;
  wire[7:0] T862;
  wire[2:0] T863;
  wire[1:0] T864;
  wire T865;
  wire[5:0] T866;
  wire[5:0] T867;
  wire[5:0] tgtPagesOH_33;
  wire[7:0] T868;
  wire[2:0] T869;
  wire T870;
  wire[5:0] T871;
  wire[5:0] T872;
  wire[5:0] tgtPagesOH_34;
  wire[7:0] T873;
  wire[2:0] T874;
  wire[3:0] T875;
  wire[1:0] T876;
  wire T877;
  wire[5:0] T878;
  wire[5:0] T879;
  wire[5:0] tgtPagesOH_35;
  wire[7:0] T880;
  wire[2:0] T881;
  wire T882;
  wire[5:0] T883;
  wire[5:0] T884;
  wire[5:0] tgtPagesOH_36;
  wire[7:0] T885;
  wire[2:0] T886;
  wire[1:0] T887;
  wire T888;
  wire[5:0] T889;
  wire[5:0] T890;
  wire[5:0] tgtPagesOH_37;
  wire[7:0] T891;
  wire[2:0] T892;
  wire T893;
  wire[5:0] T894;
  wire[5:0] T895;
  wire[5:0] tgtPagesOH_38;
  wire[7:0] T896;
  wire[2:0] T897;
  wire[7:0] T898;
  wire[3:0] T899;
  wire[1:0] T900;
  wire T901;
  wire[5:0] T902;
  wire[5:0] T903;
  wire[5:0] tgtPagesOH_39;
  wire[7:0] T904;
  wire[2:0] T905;
  wire T906;
  wire[5:0] T907;
  wire[5:0] T908;
  wire[5:0] tgtPagesOH_40;
  wire[7:0] T909;
  wire[2:0] T910;
  wire[1:0] T911;
  wire T912;
  wire[5:0] T913;
  wire[5:0] T914;
  wire[5:0] tgtPagesOH_41;
  wire[7:0] T915;
  wire[2:0] T916;
  wire T917;
  wire[5:0] T918;
  wire[5:0] T919;
  wire[5:0] tgtPagesOH_42;
  wire[7:0] T920;
  wire[2:0] T921;
  wire[3:0] T922;
  wire[1:0] T923;
  wire T924;
  wire[5:0] T925;
  wire[5:0] T926;
  wire[5:0] tgtPagesOH_43;
  wire[7:0] T927;
  wire[2:0] T928;
  wire T929;
  wire[5:0] T930;
  wire[5:0] T931;
  wire[5:0] tgtPagesOH_44;
  wire[7:0] T932;
  wire[2:0] T933;
  wire[1:0] T934;
  wire T935;
  wire[5:0] T936;
  wire[5:0] T937;
  wire[5:0] tgtPagesOH_45;
  wire[7:0] T938;
  wire[2:0] T939;
  wire T940;
  wire[5:0] T941;
  wire[5:0] T942;
  wire[5:0] tgtPagesOH_46;
  wire[7:0] T943;
  wire[2:0] T944;
  wire[14:0] T945;
  wire[7:0] T946;
  wire[3:0] T947;
  wire[1:0] T948;
  wire T949;
  wire[5:0] T950;
  wire[5:0] T951;
  wire[5:0] tgtPagesOH_47;
  wire[7:0] T952;
  wire[2:0] T953;
  wire T954;
  wire[5:0] T955;
  wire[5:0] T956;
  wire[5:0] tgtPagesOH_48;
  wire[7:0] T957;
  wire[2:0] T958;
  wire[1:0] T959;
  wire T960;
  wire[5:0] T961;
  wire[5:0] T962;
  wire[5:0] tgtPagesOH_49;
  wire[7:0] T963;
  wire[2:0] T964;
  wire T965;
  wire[5:0] T966;
  wire[5:0] T967;
  wire[5:0] tgtPagesOH_50;
  wire[7:0] T968;
  wire[2:0] T969;
  wire[3:0] T970;
  wire[1:0] T971;
  wire T972;
  wire[5:0] T973;
  wire[5:0] T974;
  wire[5:0] tgtPagesOH_51;
  wire[7:0] T975;
  wire[2:0] T976;
  wire T977;
  wire[5:0] T978;
  wire[5:0] T979;
  wire[5:0] tgtPagesOH_52;
  wire[7:0] T980;
  wire[2:0] T981;
  wire[1:0] T982;
  wire T983;
  wire[5:0] T984;
  wire[5:0] T985;
  wire[5:0] tgtPagesOH_53;
  wire[7:0] T986;
  wire[2:0] T987;
  wire T988;
  wire[5:0] T989;
  wire[5:0] T990;
  wire[5:0] tgtPagesOH_54;
  wire[7:0] T991;
  wire[2:0] T992;
  wire[6:0] T993;
  wire[3:0] T994;
  wire[1:0] T995;
  wire T996;
  wire[5:0] T997;
  wire[5:0] T998;
  wire[5:0] tgtPagesOH_55;
  wire[7:0] T999;
  wire[2:0] T1000;
  wire T1001;
  wire[5:0] T1002;
  wire[5:0] T1003;
  wire[5:0] tgtPagesOH_56;
  wire[7:0] T1004;
  wire[2:0] T1005;
  wire[1:0] T1006;
  wire T1007;
  wire[5:0] T1008;
  wire[5:0] T1009;
  wire[5:0] tgtPagesOH_57;
  wire[7:0] T1010;
  wire[2:0] T1011;
  wire T1012;
  wire[5:0] T1013;
  wire[5:0] T1014;
  wire[5:0] tgtPagesOH_58;
  wire[7:0] T1015;
  wire[2:0] T1016;
  wire[2:0] T1017;
  wire[1:0] T1018;
  wire T1019;
  wire[5:0] T1020;
  wire[5:0] T1021;
  wire[5:0] tgtPagesOH_59;
  wire[7:0] T1022;
  wire[2:0] T1023;
  wire T1024;
  wire[5:0] T1025;
  wire[5:0] T1026;
  wire[5:0] tgtPagesOH_60;
  wire[7:0] T1027;
  wire[2:0] T1028;
  wire T1029;
  wire[5:0] T1030;
  wire[5:0] T1031;
  wire[5:0] tgtPagesOH_61;
  wire[7:0] T1032;
  wire[2:0] T1033;
  wire T1034;
  wire T1035;
  reg  isJump_60;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  reg  isJump_59;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire T1046;
  wire T1047;
  reg  isJump_58;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire T1053;
  reg  isJump_57;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  reg  isJump_56;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  reg  isJump_55;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire T1071;
  reg  isJump_54;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  reg  isJump_53;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  reg  isJump_52;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  reg  isJump_51;
  wire T1090;
  wire T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  reg  isJump_50;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  reg  isJump_49;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  reg  isJump_48;
  wire T1108;
  wire T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  reg  isJump_47;
  wire T1114;
  wire T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  reg  isJump_46;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire T1125;
  reg  isJump_45;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  reg  isJump_44;
  wire T1132;
  wire T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  reg  isJump_43;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  reg  isJump_42;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire T1149;
  reg  isJump_41;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  reg  isJump_40;
  wire T1156;
  wire T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  reg  isJump_39;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  reg  isJump_38;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  reg  isJump_37;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  reg  isJump_36;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire T1185;
  reg  isJump_35;
  wire T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire T1191;
  reg  isJump_34;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  reg  isJump_33;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  reg  isJump_32;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire T1209;
  reg  isJump_31;
  wire T1210;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  reg  isJump_30;
  wire T1216;
  wire T1217;
  wire T1218;
  wire T1219;
  wire T1220;
  wire T1221;
  reg  isJump_29;
  wire T1222;
  wire T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  reg  isJump_28;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  reg  isJump_27;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  reg  isJump_26;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  reg  isJump_25;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  reg  isJump_24;
  wire T1252;
  wire T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire T1257;
  reg  isJump_23;
  wire T1258;
  wire T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  reg  isJump_22;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire T1268;
  wire T1269;
  reg  isJump_21;
  wire T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  reg  isJump_20;
  wire T1276;
  wire T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  reg  isJump_19;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  reg  isJump_18;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire T1292;
  wire T1293;
  reg  isJump_17;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  reg  isJump_16;
  wire T1300;
  wire T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  reg  isJump_15;
  wire T1306;
  wire T1307;
  wire T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  reg  isJump_14;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  reg  isJump_13;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  reg  isJump_12;
  wire T1324;
  wire T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  reg  isJump_11;
  wire T1330;
  wire T1331;
  wire T1332;
  wire T1333;
  wire T1334;
  wire T1335;
  reg  isJump_10;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  reg  isJump_9;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  reg  isJump_8;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire T1353;
  reg  isJump_7;
  wire T1354;
  wire T1355;
  wire T1356;
  wire T1357;
  wire T1358;
  wire T1359;
  reg  isJump_6;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire T1364;
  wire T1365;
  reg  isJump_5;
  wire T1366;
  wire T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  reg  isJump_4;
  wire T1372;
  wire T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  reg  isJump_3;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  reg  isJump_2;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  reg  isJump_1;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  reg  isJump_0;
  wire T1395;
  wire T1396;
  wire T1397;
  wire T1398;
  wire T1399;
  wire[6:0] T1400;
  wire[5:0] T1401;
  wire T1402;
  wire[6:0] T1403;
  wire[6:0] T1404;
  wire[5:0] T2321;
  wire[4:0] T2322;
  wire[3:0] T2323;
  wire[2:0] T2324;
  wire[1:0] T2325;
  wire T2326;
  wire[1:0] T2327;
  wire[1:0] T2328;
  wire[3:0] T2329;
  wire[3:0] T2330;
  wire[7:0] T2331;
  wire[7:0] T2332;
  wire[15:0] T2333;
  wire[15:0] T2334;
  wire[31:0] T2335;
  wire[31:0] T2336;
  wire[29:0] T2337;
  wire[15:0] T2338;
  wire[7:0] T2339;
  wire[3:0] T2340;
  wire[1:0] T2341;
  wire T2342;
  wire T2343;
  wire T2344;
  wire T2345;
  wire T2346;
  wire[38:0] T1406;
  wire[38:0] T1407;
  wire[38:0] T1408;
  wire[11:0] T1409;
  wire[11:0] T1410;
  wire[11:0] T1411;
  reg [11:0] tgts [61:0];
  wire[11:0] T1412;
  wire[11:0] T2347;
  wire T1413;
  wire T1414;
  wire T1415;
  wire[11:0] T1416;
  wire[11:0] T1417;
  wire[11:0] T1418;
  wire T1419;
  wire[11:0] T1420;
  wire[11:0] T1421;
  wire[11:0] T1422;
  wire T1423;
  wire[11:0] T1424;
  wire[11:0] T1425;
  wire[11:0] T1426;
  wire T1427;
  wire[11:0] T1428;
  wire[11:0] T1429;
  wire[11:0] T1430;
  wire T1431;
  wire[11:0] T1432;
  wire[11:0] T1433;
  wire[11:0] T1434;
  wire T1435;
  wire[11:0] T1436;
  wire[11:0] T1437;
  wire[11:0] T1438;
  wire T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[11:0] T1442;
  wire T1443;
  wire[11:0] T1444;
  wire[11:0] T1445;
  wire[11:0] T1446;
  wire T1447;
  wire[11:0] T1448;
  wire[11:0] T1449;
  wire[11:0] T1450;
  wire T1451;
  wire[11:0] T1452;
  wire[11:0] T1453;
  wire[11:0] T1454;
  wire T1455;
  wire[11:0] T1456;
  wire[11:0] T1457;
  wire[11:0] T1458;
  wire T1459;
  wire[11:0] T1460;
  wire[11:0] T1461;
  wire[11:0] T1462;
  wire T1463;
  wire[11:0] T1464;
  wire[11:0] T1465;
  wire[11:0] T1466;
  wire T1467;
  wire[11:0] T1468;
  wire[11:0] T1469;
  wire[11:0] T1470;
  wire T1471;
  wire[11:0] T1472;
  wire[11:0] T1473;
  wire[11:0] T1474;
  wire T1475;
  wire[11:0] T1476;
  wire[11:0] T1477;
  wire[11:0] T1478;
  wire T1479;
  wire[11:0] T1480;
  wire[11:0] T1481;
  wire[11:0] T1482;
  wire T1483;
  wire[11:0] T1484;
  wire[11:0] T1485;
  wire[11:0] T1486;
  wire T1487;
  wire[11:0] T1488;
  wire[11:0] T1489;
  wire[11:0] T1490;
  wire T1491;
  wire[11:0] T1492;
  wire[11:0] T1493;
  wire[11:0] T1494;
  wire T1495;
  wire[11:0] T1496;
  wire[11:0] T1497;
  wire[11:0] T1498;
  wire T1499;
  wire[11:0] T1500;
  wire[11:0] T1501;
  wire[11:0] T1502;
  wire T1503;
  wire[11:0] T1504;
  wire[11:0] T1505;
  wire[11:0] T1506;
  wire T1507;
  wire[11:0] T1508;
  wire[11:0] T1509;
  wire[11:0] T1510;
  wire T1511;
  wire[11:0] T1512;
  wire[11:0] T1513;
  wire[11:0] T1514;
  wire T1515;
  wire[11:0] T1516;
  wire[11:0] T1517;
  wire[11:0] T1518;
  wire T1519;
  wire[11:0] T1520;
  wire[11:0] T1521;
  wire[11:0] T1522;
  wire T1523;
  wire[11:0] T1524;
  wire[11:0] T1525;
  wire[11:0] T1526;
  wire T1527;
  wire[11:0] T1528;
  wire[11:0] T1529;
  wire[11:0] T1530;
  wire T1531;
  wire[11:0] T1532;
  wire[11:0] T1533;
  wire[11:0] T1534;
  wire T1535;
  wire[11:0] T1536;
  wire[11:0] T1537;
  wire[11:0] T1538;
  wire T1539;
  wire[11:0] T1540;
  wire[11:0] T1541;
  wire[11:0] T1542;
  wire T1543;
  wire[11:0] T1544;
  wire[11:0] T1545;
  wire[11:0] T1546;
  wire T1547;
  wire[11:0] T1548;
  wire[11:0] T1549;
  wire[11:0] T1550;
  wire T1551;
  wire[11:0] T1552;
  wire[11:0] T1553;
  wire[11:0] T1554;
  wire T1555;
  wire[11:0] T1556;
  wire[11:0] T1557;
  wire[11:0] T1558;
  wire T1559;
  wire[11:0] T1560;
  wire[11:0] T1561;
  wire[11:0] T1562;
  wire T1563;
  wire[11:0] T1564;
  wire[11:0] T1565;
  wire[11:0] T1566;
  wire T1567;
  wire[11:0] T1568;
  wire[11:0] T1569;
  wire[11:0] T1570;
  wire T1571;
  wire[11:0] T1572;
  wire[11:0] T1573;
  wire[11:0] T1574;
  wire T1575;
  wire[11:0] T1576;
  wire[11:0] T1577;
  wire[11:0] T1578;
  wire T1579;
  wire[11:0] T1580;
  wire[11:0] T1581;
  wire[11:0] T1582;
  wire T1583;
  wire[11:0] T1584;
  wire[11:0] T1585;
  wire[11:0] T1586;
  wire T1587;
  wire[11:0] T1588;
  wire[11:0] T1589;
  wire[11:0] T1590;
  wire T1591;
  wire[11:0] T1592;
  wire[11:0] T1593;
  wire[11:0] T1594;
  wire T1595;
  wire[11:0] T1596;
  wire[11:0] T1597;
  wire[11:0] T1598;
  wire T1599;
  wire[11:0] T1600;
  wire[11:0] T1601;
  wire[11:0] T1602;
  wire T1603;
  wire[11:0] T1604;
  wire[11:0] T1605;
  wire[11:0] T1606;
  wire T1607;
  wire[11:0] T1608;
  wire[11:0] T1609;
  wire[11:0] T1610;
  wire T1611;
  wire[11:0] T1612;
  wire[11:0] T1613;
  wire[11:0] T1614;
  wire T1615;
  wire[11:0] T1616;
  wire[11:0] T1617;
  wire[11:0] T1618;
  wire T1619;
  wire[11:0] T1620;
  wire[11:0] T1621;
  wire[11:0] T1622;
  wire T1623;
  wire[11:0] T1624;
  wire[11:0] T1625;
  wire[11:0] T1626;
  wire T1627;
  wire[11:0] T1628;
  wire[11:0] T1629;
  wire[11:0] T1630;
  wire T1631;
  wire[11:0] T1632;
  wire[11:0] T1633;
  wire[11:0] T1634;
  wire T1635;
  wire[11:0] T1636;
  wire[11:0] T1637;
  wire[11:0] T1638;
  wire T1639;
  wire[11:0] T1640;
  wire[11:0] T1641;
  wire[11:0] T1642;
  wire T1643;
  wire[11:0] T1644;
  wire[11:0] T1645;
  wire[11:0] T1646;
  wire T1647;
  wire[11:0] T1648;
  wire[11:0] T1649;
  wire[11:0] T1650;
  wire T1651;
  wire[11:0] T1652;
  wire[11:0] T1653;
  wire[11:0] T1654;
  wire T1655;
  wire[11:0] T1656;
  wire[11:0] T1657;
  wire T1658;
  wire[26:0] T1659;
  wire[26:0] T1660;
  wire[26:0] T1661;
  wire T1662;
  wire[5:0] T1663;
  wire[5:0] T1664;
  wire T1665;
  wire[5:0] T1666;
  wire[5:0] T1667;
  wire T1668;
  wire[5:0] T1669;
  wire[5:0] T1670;
  wire T1671;
  wire[5:0] T1672;
  wire[5:0] T1673;
  wire T1674;
  wire[5:0] T1675;
  wire[5:0] T1676;
  wire T1677;
  wire[5:0] T1678;
  wire[5:0] T1679;
  wire T1680;
  wire[5:0] T1681;
  wire[5:0] T1682;
  wire T1683;
  wire[5:0] T1684;
  wire[5:0] T1685;
  wire T1686;
  wire[5:0] T1687;
  wire[5:0] T1688;
  wire T1689;
  wire[5:0] T1690;
  wire[5:0] T1691;
  wire T1692;
  wire[5:0] T1693;
  wire[5:0] T1694;
  wire T1695;
  wire[5:0] T1696;
  wire[5:0] T1697;
  wire T1698;
  wire[5:0] T1699;
  wire[5:0] T1700;
  wire T1701;
  wire[5:0] T1702;
  wire[5:0] T1703;
  wire T1704;
  wire[5:0] T1705;
  wire[5:0] T1706;
  wire T1707;
  wire[5:0] T1708;
  wire[5:0] T1709;
  wire T1710;
  wire[5:0] T1711;
  wire[5:0] T1712;
  wire T1713;
  wire[5:0] T1714;
  wire[5:0] T1715;
  wire T1716;
  wire[5:0] T1717;
  wire[5:0] T1718;
  wire T1719;
  wire[5:0] T1720;
  wire[5:0] T1721;
  wire T1722;
  wire[5:0] T1723;
  wire[5:0] T1724;
  wire T1725;
  wire[5:0] T1726;
  wire[5:0] T1727;
  wire T1728;
  wire[5:0] T1729;
  wire[5:0] T1730;
  wire T1731;
  wire[5:0] T1732;
  wire[5:0] T1733;
  wire T1734;
  wire[5:0] T1735;
  wire[5:0] T1736;
  wire T1737;
  wire[5:0] T1738;
  wire[5:0] T1739;
  wire T1740;
  wire[5:0] T1741;
  wire[5:0] T1742;
  wire T1743;
  wire[5:0] T1744;
  wire[5:0] T1745;
  wire T1746;
  wire[5:0] T1747;
  wire[5:0] T1748;
  wire T1749;
  wire[5:0] T1750;
  wire[5:0] T1751;
  wire T1752;
  wire[5:0] T1753;
  wire[5:0] T1754;
  wire T1755;
  wire[5:0] T1756;
  wire[5:0] T1757;
  wire T1758;
  wire[5:0] T1759;
  wire[5:0] T1760;
  wire T1761;
  wire[5:0] T1762;
  wire[5:0] T1763;
  wire T1764;
  wire[5:0] T1765;
  wire[5:0] T1766;
  wire T1767;
  wire[5:0] T1768;
  wire[5:0] T1769;
  wire T1770;
  wire[5:0] T1771;
  wire[5:0] T1772;
  wire T1773;
  wire[5:0] T1774;
  wire[5:0] T1775;
  wire T1776;
  wire[5:0] T1777;
  wire[5:0] T1778;
  wire T1779;
  wire[5:0] T1780;
  wire[5:0] T1781;
  wire T1782;
  wire[5:0] T1783;
  wire[5:0] T1784;
  wire T1785;
  wire[5:0] T1786;
  wire[5:0] T1787;
  wire T1788;
  wire[5:0] T1789;
  wire[5:0] T1790;
  wire T1791;
  wire[5:0] T1792;
  wire[5:0] T1793;
  wire T1794;
  wire[5:0] T1795;
  wire[5:0] T1796;
  wire T1797;
  wire[5:0] T1798;
  wire[5:0] T1799;
  wire T1800;
  wire[5:0] T1801;
  wire[5:0] T1802;
  wire T1803;
  wire[5:0] T1804;
  wire[5:0] T1805;
  wire T1806;
  wire[5:0] T1807;
  wire[5:0] T1808;
  wire T1809;
  wire[5:0] T1810;
  wire[5:0] T1811;
  wire T1812;
  wire[5:0] T1813;
  wire[5:0] T1814;
  wire T1815;
  wire[5:0] T1816;
  wire[5:0] T1817;
  wire T1818;
  wire[5:0] T1819;
  wire[5:0] T1820;
  wire T1821;
  wire[5:0] T1822;
  wire[5:0] T1823;
  wire T1824;
  wire[5:0] T1825;
  wire[5:0] T1826;
  wire T1827;
  wire[5:0] T1828;
  wire[5:0] T1829;
  wire T1830;
  wire[5:0] T1831;
  wire[5:0] T1832;
  wire T1833;
  wire[5:0] T1834;
  wire[5:0] T1835;
  wire T1836;
  wire[5:0] T1837;
  wire[5:0] T1838;
  wire T1839;
  wire[5:0] T1840;
  wire[5:0] T1841;
  wire T1842;
  wire[5:0] T1843;
  wire[5:0] T1844;
  wire T1845;
  wire[5:0] T1846;
  wire T1847;
  wire[26:0] T1848;
  wire[26:0] T1849;
  wire[26:0] T1850;
  wire T1851;
  wire[26:0] T1852;
  wire[26:0] T1853;
  wire[26:0] T1854;
  wire T1855;
  wire[26:0] T1856;
  wire[26:0] T1857;
  wire[26:0] T1858;
  wire T1859;
  wire[26:0] T1860;
  wire[26:0] T1861;
  wire[26:0] T1862;
  wire T1863;
  wire[26:0] T1864;
  wire[26:0] T1865;
  wire T1866;
  wire[38:0] T1867;
  reg [38:0] R1868;
  wire[38:0] T1869;
  wire T1870;
  wire T1871;
  wire[1:0] T1872;
  wire T1873;
  wire T1874;
  reg  R1875;
  wire T2348;
  wire T1876;
  wire T1877;
  wire T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  reg [1:0] R1882;
  wire[1:0] T2349;
  wire[1:0] T1883;
  wire[1:0] T1884;
  wire[1:0] T1885;
  wire[1:0] T1886;
  wire T1887;
  wire T1888;
  wire[1:0] T1889;
  wire T1890;
  wire T1891;
  wire T1892;
  wire T1893;
  wire T1894;
  reg [38:0] R1895;
  wire[38:0] T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire T1900;
  wire T1901;
  wire T1902;
  reg  useRAS_61;
  wire T1903;
  reg  R1904;
  wire T1905;
  wire T1906;
  wire T1907;
  wire[63:0] T1908;
  wire[5:0] T1909;
  wire T1910;
  wire T1911;
  wire T1912;
  reg  useRAS_60;
  wire T1913;
  wire T1914;
  wire T1915;
  wire T1916;
  wire T1917;
  wire T1918;
  reg  useRAS_59;
  wire T1919;
  wire T1920;
  wire T1921;
  wire T1922;
  wire T1923;
  wire T1924;
  reg  useRAS_58;
  wire T1925;
  wire T1926;
  wire T1927;
  wire T1928;
  wire T1929;
  wire T1930;
  reg  useRAS_57;
  wire T1931;
  wire T1932;
  wire T1933;
  wire T1934;
  wire T1935;
  wire T1936;
  reg  useRAS_56;
  wire T1937;
  wire T1938;
  wire T1939;
  wire T1940;
  wire T1941;
  wire T1942;
  reg  useRAS_55;
  wire T1943;
  wire T1944;
  wire T1945;
  wire T1946;
  wire T1947;
  wire T1948;
  reg  useRAS_54;
  wire T1949;
  wire T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire T1954;
  reg  useRAS_53;
  wire T1955;
  wire T1956;
  wire T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  reg  useRAS_52;
  wire T1961;
  wire T1962;
  wire T1963;
  wire T1964;
  wire T1965;
  wire T1966;
  reg  useRAS_51;
  wire T1967;
  wire T1968;
  wire T1969;
  wire T1970;
  wire T1971;
  wire T1972;
  reg  useRAS_50;
  wire T1973;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  reg  useRAS_49;
  wire T1979;
  wire T1980;
  wire T1981;
  wire T1982;
  wire T1983;
  wire T1984;
  reg  useRAS_48;
  wire T1985;
  wire T1986;
  wire T1987;
  wire T1988;
  wire T1989;
  wire T1990;
  reg  useRAS_47;
  wire T1991;
  wire T1992;
  wire T1993;
  wire T1994;
  wire T1995;
  wire T1996;
  reg  useRAS_46;
  wire T1997;
  wire T1998;
  wire T1999;
  wire T2000;
  wire T2001;
  wire T2002;
  reg  useRAS_45;
  wire T2003;
  wire T2004;
  wire T2005;
  wire T2006;
  wire T2007;
  wire T2008;
  reg  useRAS_44;
  wire T2009;
  wire T2010;
  wire T2011;
  wire T2012;
  wire T2013;
  wire T2014;
  reg  useRAS_43;
  wire T2015;
  wire T2016;
  wire T2017;
  wire T2018;
  wire T2019;
  wire T2020;
  reg  useRAS_42;
  wire T2021;
  wire T2022;
  wire T2023;
  wire T2024;
  wire T2025;
  wire T2026;
  reg  useRAS_41;
  wire T2027;
  wire T2028;
  wire T2029;
  wire T2030;
  wire T2031;
  wire T2032;
  reg  useRAS_40;
  wire T2033;
  wire T2034;
  wire T2035;
  wire T2036;
  wire T2037;
  wire T2038;
  reg  useRAS_39;
  wire T2039;
  wire T2040;
  wire T2041;
  wire T2042;
  wire T2043;
  wire T2044;
  reg  useRAS_38;
  wire T2045;
  wire T2046;
  wire T2047;
  wire T2048;
  wire T2049;
  wire T2050;
  reg  useRAS_37;
  wire T2051;
  wire T2052;
  wire T2053;
  wire T2054;
  wire T2055;
  wire T2056;
  reg  useRAS_36;
  wire T2057;
  wire T2058;
  wire T2059;
  wire T2060;
  wire T2061;
  wire T2062;
  reg  useRAS_35;
  wire T2063;
  wire T2064;
  wire T2065;
  wire T2066;
  wire T2067;
  wire T2068;
  reg  useRAS_34;
  wire T2069;
  wire T2070;
  wire T2071;
  wire T2072;
  wire T2073;
  wire T2074;
  reg  useRAS_33;
  wire T2075;
  wire T2076;
  wire T2077;
  wire T2078;
  wire T2079;
  wire T2080;
  reg  useRAS_32;
  wire T2081;
  wire T2082;
  wire T2083;
  wire T2084;
  wire T2085;
  wire T2086;
  reg  useRAS_31;
  wire T2087;
  wire T2088;
  wire T2089;
  wire T2090;
  wire T2091;
  wire T2092;
  reg  useRAS_30;
  wire T2093;
  wire T2094;
  wire T2095;
  wire T2096;
  wire T2097;
  wire T2098;
  reg  useRAS_29;
  wire T2099;
  wire T2100;
  wire T2101;
  wire T2102;
  wire T2103;
  wire T2104;
  reg  useRAS_28;
  wire T2105;
  wire T2106;
  wire T2107;
  wire T2108;
  wire T2109;
  wire T2110;
  reg  useRAS_27;
  wire T2111;
  wire T2112;
  wire T2113;
  wire T2114;
  wire T2115;
  wire T2116;
  reg  useRAS_26;
  wire T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire T2121;
  wire T2122;
  reg  useRAS_25;
  wire T2123;
  wire T2124;
  wire T2125;
  wire T2126;
  wire T2127;
  wire T2128;
  reg  useRAS_24;
  wire T2129;
  wire T2130;
  wire T2131;
  wire T2132;
  wire T2133;
  wire T2134;
  reg  useRAS_23;
  wire T2135;
  wire T2136;
  wire T2137;
  wire T2138;
  wire T2139;
  wire T2140;
  reg  useRAS_22;
  wire T2141;
  wire T2142;
  wire T2143;
  wire T2144;
  wire T2145;
  wire T2146;
  reg  useRAS_21;
  wire T2147;
  wire T2148;
  wire T2149;
  wire T2150;
  wire T2151;
  wire T2152;
  reg  useRAS_20;
  wire T2153;
  wire T2154;
  wire T2155;
  wire T2156;
  wire T2157;
  wire T2158;
  reg  useRAS_19;
  wire T2159;
  wire T2160;
  wire T2161;
  wire T2162;
  wire T2163;
  wire T2164;
  reg  useRAS_18;
  wire T2165;
  wire T2166;
  wire T2167;
  wire T2168;
  wire T2169;
  wire T2170;
  reg  useRAS_17;
  wire T2171;
  wire T2172;
  wire T2173;
  wire T2174;
  wire T2175;
  wire T2176;
  reg  useRAS_16;
  wire T2177;
  wire T2178;
  wire T2179;
  wire T2180;
  wire T2181;
  wire T2182;
  reg  useRAS_15;
  wire T2183;
  wire T2184;
  wire T2185;
  wire T2186;
  wire T2187;
  wire T2188;
  reg  useRAS_14;
  wire T2189;
  wire T2190;
  wire T2191;
  wire T2192;
  wire T2193;
  wire T2194;
  reg  useRAS_13;
  wire T2195;
  wire T2196;
  wire T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  reg  useRAS_12;
  wire T2201;
  wire T2202;
  wire T2203;
  wire T2204;
  wire T2205;
  wire T2206;
  reg  useRAS_11;
  wire T2207;
  wire T2208;
  wire T2209;
  wire T2210;
  wire T2211;
  wire T2212;
  reg  useRAS_10;
  wire T2213;
  wire T2214;
  wire T2215;
  wire T2216;
  wire T2217;
  wire T2218;
  reg  useRAS_9;
  wire T2219;
  wire T2220;
  wire T2221;
  wire T2222;
  wire T2223;
  wire T2224;
  reg  useRAS_8;
  wire T2225;
  wire T2226;
  wire T2227;
  wire T2228;
  wire T2229;
  wire T2230;
  reg  useRAS_7;
  wire T2231;
  wire T2232;
  wire T2233;
  wire T2234;
  wire T2235;
  wire T2236;
  reg  useRAS_6;
  wire T2237;
  wire T2238;
  wire T2239;
  wire T2240;
  wire T2241;
  wire T2242;
  reg  useRAS_5;
  wire T2243;
  wire T2244;
  wire T2245;
  wire T2246;
  wire T2247;
  wire T2248;
  reg  useRAS_4;
  wire T2249;
  wire T2250;
  wire T2251;
  wire T2252;
  wire T2253;
  wire T2254;
  reg  useRAS_3;
  wire T2255;
  wire T2256;
  wire T2257;
  wire T2258;
  wire T2259;
  wire T2260;
  reg  useRAS_2;
  wire T2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire T2265;
  wire T2266;
  reg  useRAS_1;
  wire T2267;
  wire T2268;
  wire T2269;
  wire T2270;
  wire T2271;
  reg  useRAS_0;
  wire T2272;
  wire T2273;
  wire T2274;
  wire T2275;
  wire T2276;
  wire T2277;
  wire T2278;
  wire T2279;
  reg [0:0] brIdx [61:0];
  wire T2280;
  wire T2281;
  wire T2282;
  wire T2283;
  wire T2284;
  wire T2285;
  wire T2286;
  wire T2287;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {2{$random}};
    R7 = {1{$random}};
    for (initvar = 0; initvar < 128; initvar = initvar+1)
      T10[initvar] = {1{$random}};
    R25 = {1{$random}};
    isJump_61 = {1{$random}};
    R36 = {1{$random}};
    nextRepl = {1{$random}};
    R49 = {1{$random}};
    updateHit = {1{$random}};
    pageValid = {1{$random}};
    R70 = {1{$random}};
    R82 = {2{$random}};
    for (initvar = 0; initvar < 6; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {2{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    isJump_60 = {1{$random}};
    isJump_59 = {1{$random}};
    isJump_58 = {1{$random}};
    isJump_57 = {1{$random}};
    isJump_56 = {1{$random}};
    isJump_55 = {1{$random}};
    isJump_54 = {1{$random}};
    isJump_53 = {1{$random}};
    isJump_52 = {1{$random}};
    isJump_51 = {1{$random}};
    isJump_50 = {1{$random}};
    isJump_49 = {1{$random}};
    isJump_48 = {1{$random}};
    isJump_47 = {1{$random}};
    isJump_46 = {1{$random}};
    isJump_45 = {1{$random}};
    isJump_44 = {1{$random}};
    isJump_43 = {1{$random}};
    isJump_42 = {1{$random}};
    isJump_41 = {1{$random}};
    isJump_40 = {1{$random}};
    isJump_39 = {1{$random}};
    isJump_38 = {1{$random}};
    isJump_37 = {1{$random}};
    isJump_36 = {1{$random}};
    isJump_35 = {1{$random}};
    isJump_34 = {1{$random}};
    isJump_33 = {1{$random}};
    isJump_32 = {1{$random}};
    isJump_31 = {1{$random}};
    isJump_30 = {1{$random}};
    isJump_29 = {1{$random}};
    isJump_28 = {1{$random}};
    isJump_27 = {1{$random}};
    isJump_26 = {1{$random}};
    isJump_25 = {1{$random}};
    isJump_24 = {1{$random}};
    isJump_23 = {1{$random}};
    isJump_22 = {1{$random}};
    isJump_21 = {1{$random}};
    isJump_20 = {1{$random}};
    isJump_19 = {1{$random}};
    isJump_18 = {1{$random}};
    isJump_17 = {1{$random}};
    isJump_16 = {1{$random}};
    isJump_15 = {1{$random}};
    isJump_14 = {1{$random}};
    isJump_13 = {1{$random}};
    isJump_12 = {1{$random}};
    isJump_11 = {1{$random}};
    isJump_10 = {1{$random}};
    isJump_9 = {1{$random}};
    isJump_8 = {1{$random}};
    isJump_7 = {1{$random}};
    isJump_6 = {1{$random}};
    isJump_5 = {1{$random}};
    isJump_4 = {1{$random}};
    isJump_3 = {1{$random}};
    isJump_2 = {1{$random}};
    isJump_1 = {1{$random}};
    isJump_0 = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R1868 = {2{$random}};
    R1875 = {1{$random}};
    R1882 = {1{$random}};
    R1895 = {2{$random}};
    useRAS_61 = {1{$random}};
    R1904 = {1{$random}};
    useRAS_60 = {1{$random}};
    useRAS_59 = {1{$random}};
    useRAS_58 = {1{$random}};
    useRAS_57 = {1{$random}};
    useRAS_56 = {1{$random}};
    useRAS_55 = {1{$random}};
    useRAS_54 = {1{$random}};
    useRAS_53 = {1{$random}};
    useRAS_52 = {1{$random}};
    useRAS_51 = {1{$random}};
    useRAS_50 = {1{$random}};
    useRAS_49 = {1{$random}};
    useRAS_48 = {1{$random}};
    useRAS_47 = {1{$random}};
    useRAS_46 = {1{$random}};
    useRAS_45 = {1{$random}};
    useRAS_44 = {1{$random}};
    useRAS_43 = {1{$random}};
    useRAS_42 = {1{$random}};
    useRAS_41 = {1{$random}};
    useRAS_40 = {1{$random}};
    useRAS_39 = {1{$random}};
    useRAS_38 = {1{$random}};
    useRAS_37 = {1{$random}};
    useRAS_36 = {1{$random}};
    useRAS_35 = {1{$random}};
    useRAS_34 = {1{$random}};
    useRAS_33 = {1{$random}};
    useRAS_32 = {1{$random}};
    useRAS_31 = {1{$random}};
    useRAS_30 = {1{$random}};
    useRAS_29 = {1{$random}};
    useRAS_28 = {1{$random}};
    useRAS_27 = {1{$random}};
    useRAS_26 = {1{$random}};
    useRAS_25 = {1{$random}};
    useRAS_24 = {1{$random}};
    useRAS_23 = {1{$random}};
    useRAS_22 = {1{$random}};
    useRAS_21 = {1{$random}};
    useRAS_20 = {1{$random}};
    useRAS_19 = {1{$random}};
    useRAS_18 = {1{$random}};
    useRAS_17 = {1{$random}};
    useRAS_16 = {1{$random}};
    useRAS_15 = {1{$random}};
    useRAS_14 = {1{$random}};
    useRAS_13 = {1{$random}};
    useRAS_12 = {1{$random}};
    useRAS_11 = {1{$random}};
    useRAS_10 = {1{$random}};
    useRAS_9 = {1{$random}};
    useRAS_8 = {1{$random}};
    useRAS_7 = {1{$random}};
    useRAS_6 = {1{$random}};
    useRAS_5 = {1{$random}};
    useRAS_4 = {1{$random}};
    useRAS_3 = {1{$random}};
    useRAS_2 = {1{$random}};
    useRAS_1 = {1{$random}};
    useRAS_0 = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      brIdx[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req_bits_addr == R4;
  assign T5 = io_btb_update_valid ? io_btb_update_bits_target : R4;
  assign T6 = R7 ^ 1'h1;
  assign T2288 = reset ? 1'h0 : io_btb_update_valid;
  assign io_resp_bits_bht_value = T8;
  assign T8 = T9;
  assign T9 = T10[T24];
  assign T12 = {io_bht_update_bits_taken, T13};
  assign T13 = T18 | T14;
  assign T14 = T15 & io_bht_update_bits_taken;
  assign T15 = T17 | T16;
  assign T16 = io_bht_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T17 = io_bht_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T18 = T20 & T19;
  assign T19 = io_bht_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T20 = io_bht_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T21 = io_bht_update_valid & io_bht_update_bits_prediction_valid;
  assign T22 = T23 ^ io_bht_update_bits_prediction_bits_bht_history;
  assign T23 = io_bht_update_bits_pc[4'h8:2'h2];
  assign T24 = T1403 ^ R25;
  assign T26 = T1402 ? T1400 : T27;
  assign T27 = T31 ? T28 : R25;
  assign T28 = {T30, T29};
  assign T29 = R25[3'h6:1'h1];
  assign T30 = T8[1'h0:1'h0];
  assign T31 = T1399 & T32;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T1034 | T34;
  assign T34 = T52 ? isJump_61 : 1'h0;
  assign T35 = T38 ? R36 : isJump_61;
  assign T37 = io_btb_update_valid ? io_btb_update_bits_isJump : R36;
  assign T38 = R7 & T39;
  assign T39 = T40[6'h3d:6'h3d];
  assign T40 = 1'h1 << T41;
  assign T41 = T42;
  assign T42 = updateHit ? R49 : nextRepl;
  assign T2289 = reset ? 6'h0 : T43;
  assign T43 = T47 ? T44 : nextRepl;
  assign T44 = T46 ? 6'h0 : T45;
  assign T45 = nextRepl + 6'h1;
  assign T46 = nextRepl == 6'h3d;
  assign T47 = R7 & T48;
  assign T48 = updateHit ^ 1'h1;
  assign T50 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_entry : R49;
  assign T51 = io_btb_update_valid ? io_btb_update_bits_prediction_valid : updateHit;
  assign T52 = hits[6'h3d:6'h3d];
  assign hits = T461 & T53;
  assign T53 = T54;
  assign T54 = {T307, T55};
  assign T55 = {T233, T56};
  assign T56 = {T194, T57};
  assign T57 = {T175, T58};
  assign T58 = {T166, T59};
  assign T59 = {T162, T60};
  assign T60 = T61 != 6'h0;
  assign T61 = idxPagesOH_0 & pageHit;
  assign pageHit = T138 & pageValid;
  assign T2290 = reset ? 6'h0 : T62;
  assign T62 = io_invalidate ? 6'h0 : T63;
  assign T63 = T137 ? T64 : pageValid;
  assign T64 = pageValid | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 6'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T65;
  assign T65 = T67 | T2291;
  assign T2291 = {5'h0, T66};
  assign T66 = idxPageUpdateOH[3'h5:3'h5];
  assign T67 = T68 << 1'h1;
  assign T68 = idxPageUpdateOH[3'h4:1'h0];
  assign idxPageUpdateOH = useUpdatePageHit ? updatePageHit : idxPageRepl;
  assign idxPageRepl = T2292;
  assign T2292 = T69[3'h5:1'h0];
  assign T69 = 1'h1 << R70;
  assign T2293 = reset ? 3'h0 : T71;
  assign T71 = T75 ? T72 : R70;
  assign T72 = T74 ? 3'h0 : T73;
  assign T73 = R70 + 3'h1;
  assign T74 = R70 == 3'h5;
  assign T75 = R7 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doIdxPageRepl = useUpdatePageHit ^ 1'h1;
  assign updatePageHit = T76 & pageValid;
  assign T76 = T77;
  assign T77 = {T123, T78};
  assign T78 = {T121, T79};
  assign T79 = {T119, T80};
  assign T80 = T84 == T81;
  assign T81 = R82 >> 4'hc;
  assign T83 = io_btb_update_valid ? io_btb_update_bits_pc : R82;
  assign T84 = pages[3'h0];
  assign T86 = T89 ? T88 : T87;
  assign T87 = R82 >> 4'hc;
  assign T88 = io_req_bits_addr >> 4'hc;
  assign T89 = T90 != 6'h0;
  assign T90 = idxPageUpdateOH & 6'h15;
  assign T91 = R7 & T92;
  assign T92 = T94 & T93;
  assign T93 = pageReplEn[3'h5:3'h5];
  assign T94 = T89 ? doTgtPageRepl : doIdxPageRepl;
  assign T96 = R7 & T97;
  assign T97 = T94 & T98;
  assign T98 = pageReplEn[2'h3:2'h3];
  assign T100 = R7 & T101;
  assign T101 = T94 & T102;
  assign T102 = pageReplEn[1'h1:1'h1];
  assign T104 = T89 ? T106 : T105;
  assign T105 = io_req_bits_addr >> 4'hc;
  assign T106 = R82 >> 4'hc;
  assign T107 = R7 & T108;
  assign T108 = T110 & T109;
  assign T109 = pageReplEn[3'h4:3'h4];
  assign T110 = T89 ? doIdxPageRepl : doTgtPageRepl;
  assign T112 = R7 & T113;
  assign T113 = T110 & T114;
  assign T114 = pageReplEn[2'h2:2'h2];
  assign T116 = R7 & T117;
  assign T117 = T110 & T118;
  assign T118 = pageReplEn[1'h0:1'h0];
  assign T119 = T120 == T81;
  assign T120 = pages[3'h1];
  assign T121 = T122 == T81;
  assign T122 = pages[3'h2];
  assign T123 = {T129, T124};
  assign T124 = {T127, T125};
  assign T125 = T126 == T81;
  assign T126 = pages[3'h3];
  assign T127 = T128 == T81;
  assign T128 = pages[3'h4];
  assign T129 = T130 == T81;
  assign T130 = pages[3'h5];
  assign useUpdatePageHit = updatePageHit != 6'h0;
  assign samePage = T132 == T131;
  assign T131 = io_req_bits_addr >> 4'hc;
  assign T132 = R82 >> 4'hc;
  assign doTgtPageRepl = T136 & T133;
  assign T133 = usePageHit ^ 1'h1;
  assign usePageHit = T134 != 6'h0;
  assign T134 = pageHit & T135;
  assign T135 = ~ idxPageReplEn;
  assign T136 = samePage ^ 1'h1;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 6'h0;
  assign T137 = R7 & doPageRepl;
  assign T138 = T139;
  assign T139 = {T149, T140};
  assign T140 = {T147, T141};
  assign T141 = {T145, T142};
  assign T142 = T144 == T143;
  assign T143 = io_req_bits_addr >> 4'hc;
  assign T144 = pages[3'h0];
  assign T145 = T146 == T143;
  assign T146 = pages[3'h1];
  assign T147 = T148 == T143;
  assign T148 = pages[3'h2];
  assign T149 = {T155, T150};
  assign T150 = {T153, T151};
  assign T151 = T152 == T143;
  assign T152 = pages[3'h3];
  assign T153 = T154 == T143;
  assign T154 = pages[3'h4];
  assign T155 = T156 == T143;
  assign T156 = pages[3'h5];
  assign idxPagesOH_0 = T157[3'h5:1'h0];
  assign T157 = 1'h1 << T158;
  assign T158 = idxPages[6'h0];
  assign T2294 = {T2304, T2295};
  assign T2295 = {T2303, T2296};
  assign T2296 = T2297[1'h1:1'h1];
  assign T2297 = T2302 | T2298;
  assign T2298 = T2299[1'h1:1'h0];
  assign T2299 = T2301 | T2300;
  assign T2300 = idxPageUpdateOH[2'h3:1'h0];
  assign T2301 = idxPageUpdateOH[3'h5:3'h4];
  assign T2302 = T2299[2'h3:2'h2];
  assign T2303 = T2302 != 2'h0;
  assign T2304 = T2301 != 2'h0;
  assign T160 = R7 & T161;
  assign T161 = T42 < 6'h3e;
  assign T162 = T163 != 6'h0;
  assign T163 = idxPagesOH_1 & pageHit;
  assign idxPagesOH_1 = T164[3'h5:1'h0];
  assign T164 = 1'h1 << T165;
  assign T165 = idxPages[6'h1];
  assign T166 = {T171, T167};
  assign T167 = T168 != 6'h0;
  assign T168 = idxPagesOH_2 & pageHit;
  assign idxPagesOH_2 = T169[3'h5:1'h0];
  assign T169 = 1'h1 << T170;
  assign T170 = idxPages[6'h2];
  assign T171 = T172 != 6'h0;
  assign T172 = idxPagesOH_3 & pageHit;
  assign idxPagesOH_3 = T173[3'h5:1'h0];
  assign T173 = 1'h1 << T174;
  assign T174 = idxPages[6'h3];
  assign T175 = {T185, T176};
  assign T176 = {T181, T177};
  assign T177 = T178 != 6'h0;
  assign T178 = idxPagesOH_4 & pageHit;
  assign idxPagesOH_4 = T179[3'h5:1'h0];
  assign T179 = 1'h1 << T180;
  assign T180 = idxPages[6'h4];
  assign T181 = T182 != 6'h0;
  assign T182 = idxPagesOH_5 & pageHit;
  assign idxPagesOH_5 = T183[3'h5:1'h0];
  assign T183 = 1'h1 << T184;
  assign T184 = idxPages[6'h5];
  assign T185 = {T190, T186};
  assign T186 = T187 != 6'h0;
  assign T187 = idxPagesOH_6 & pageHit;
  assign idxPagesOH_6 = T188[3'h5:1'h0];
  assign T188 = 1'h1 << T189;
  assign T189 = idxPages[6'h6];
  assign T190 = T191 != 6'h0;
  assign T191 = idxPagesOH_7 & pageHit;
  assign idxPagesOH_7 = T192[3'h5:1'h0];
  assign T192 = 1'h1 << T193;
  assign T193 = idxPages[6'h7];
  assign T194 = {T214, T195};
  assign T195 = {T205, T196};
  assign T196 = {T201, T197};
  assign T197 = T198 != 6'h0;
  assign T198 = idxPagesOH_8 & pageHit;
  assign idxPagesOH_8 = T199[3'h5:1'h0];
  assign T199 = 1'h1 << T200;
  assign T200 = idxPages[6'h8];
  assign T201 = T202 != 6'h0;
  assign T202 = idxPagesOH_9 & pageHit;
  assign idxPagesOH_9 = T203[3'h5:1'h0];
  assign T203 = 1'h1 << T204;
  assign T204 = idxPages[6'h9];
  assign T205 = {T210, T206};
  assign T206 = T207 != 6'h0;
  assign T207 = idxPagesOH_10 & pageHit;
  assign idxPagesOH_10 = T208[3'h5:1'h0];
  assign T208 = 1'h1 << T209;
  assign T209 = idxPages[6'ha];
  assign T210 = T211 != 6'h0;
  assign T211 = idxPagesOH_11 & pageHit;
  assign idxPagesOH_11 = T212[3'h5:1'h0];
  assign T212 = 1'h1 << T213;
  assign T213 = idxPages[6'hb];
  assign T214 = {T224, T215};
  assign T215 = {T220, T216};
  assign T216 = T217 != 6'h0;
  assign T217 = idxPagesOH_12 & pageHit;
  assign idxPagesOH_12 = T218[3'h5:1'h0];
  assign T218 = 1'h1 << T219;
  assign T219 = idxPages[6'hc];
  assign T220 = T221 != 6'h0;
  assign T221 = idxPagesOH_13 & pageHit;
  assign idxPagesOH_13 = T222[3'h5:1'h0];
  assign T222 = 1'h1 << T223;
  assign T223 = idxPages[6'hd];
  assign T224 = {T229, T225};
  assign T225 = T226 != 6'h0;
  assign T226 = idxPagesOH_14 & pageHit;
  assign idxPagesOH_14 = T227[3'h5:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = idxPages[6'he];
  assign T229 = T230 != 6'h0;
  assign T230 = idxPagesOH_15 & pageHit;
  assign idxPagesOH_15 = T231[3'h5:1'h0];
  assign T231 = 1'h1 << T232;
  assign T232 = idxPages[6'hf];
  assign T233 = {T273, T234};
  assign T234 = {T254, T235};
  assign T235 = {T245, T236};
  assign T236 = {T241, T237};
  assign T237 = T238 != 6'h0;
  assign T238 = idxPagesOH_16 & pageHit;
  assign idxPagesOH_16 = T239[3'h5:1'h0];
  assign T239 = 1'h1 << T240;
  assign T240 = idxPages[6'h10];
  assign T241 = T242 != 6'h0;
  assign T242 = idxPagesOH_17 & pageHit;
  assign idxPagesOH_17 = T243[3'h5:1'h0];
  assign T243 = 1'h1 << T244;
  assign T244 = idxPages[6'h11];
  assign T245 = {T250, T246};
  assign T246 = T247 != 6'h0;
  assign T247 = idxPagesOH_18 & pageHit;
  assign idxPagesOH_18 = T248[3'h5:1'h0];
  assign T248 = 1'h1 << T249;
  assign T249 = idxPages[6'h12];
  assign T250 = T251 != 6'h0;
  assign T251 = idxPagesOH_19 & pageHit;
  assign idxPagesOH_19 = T252[3'h5:1'h0];
  assign T252 = 1'h1 << T253;
  assign T253 = idxPages[6'h13];
  assign T254 = {T264, T255};
  assign T255 = {T260, T256};
  assign T256 = T257 != 6'h0;
  assign T257 = idxPagesOH_20 & pageHit;
  assign idxPagesOH_20 = T258[3'h5:1'h0];
  assign T258 = 1'h1 << T259;
  assign T259 = idxPages[6'h14];
  assign T260 = T261 != 6'h0;
  assign T261 = idxPagesOH_21 & pageHit;
  assign idxPagesOH_21 = T262[3'h5:1'h0];
  assign T262 = 1'h1 << T263;
  assign T263 = idxPages[6'h15];
  assign T264 = {T269, T265};
  assign T265 = T266 != 6'h0;
  assign T266 = idxPagesOH_22 & pageHit;
  assign idxPagesOH_22 = T267[3'h5:1'h0];
  assign T267 = 1'h1 << T268;
  assign T268 = idxPages[6'h16];
  assign T269 = T270 != 6'h0;
  assign T270 = idxPagesOH_23 & pageHit;
  assign idxPagesOH_23 = T271[3'h5:1'h0];
  assign T271 = 1'h1 << T272;
  assign T272 = idxPages[6'h17];
  assign T273 = {T293, T274};
  assign T274 = {T284, T275};
  assign T275 = {T280, T276};
  assign T276 = T277 != 6'h0;
  assign T277 = idxPagesOH_24 & pageHit;
  assign idxPagesOH_24 = T278[3'h5:1'h0];
  assign T278 = 1'h1 << T279;
  assign T279 = idxPages[6'h18];
  assign T280 = T281 != 6'h0;
  assign T281 = idxPagesOH_25 & pageHit;
  assign idxPagesOH_25 = T282[3'h5:1'h0];
  assign T282 = 1'h1 << T283;
  assign T283 = idxPages[6'h19];
  assign T284 = {T289, T285};
  assign T285 = T286 != 6'h0;
  assign T286 = idxPagesOH_26 & pageHit;
  assign idxPagesOH_26 = T287[3'h5:1'h0];
  assign T287 = 1'h1 << T288;
  assign T288 = idxPages[6'h1a];
  assign T289 = T290 != 6'h0;
  assign T290 = idxPagesOH_27 & pageHit;
  assign idxPagesOH_27 = T291[3'h5:1'h0];
  assign T291 = 1'h1 << T292;
  assign T292 = idxPages[6'h1b];
  assign T293 = {T303, T294};
  assign T294 = {T299, T295};
  assign T295 = T296 != 6'h0;
  assign T296 = idxPagesOH_28 & pageHit;
  assign idxPagesOH_28 = T297[3'h5:1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = idxPages[6'h1c];
  assign T299 = T300 != 6'h0;
  assign T300 = idxPagesOH_29 & pageHit;
  assign idxPagesOH_29 = T301[3'h5:1'h0];
  assign T301 = 1'h1 << T302;
  assign T302 = idxPages[6'h1d];
  assign T303 = T304 != 6'h0;
  assign T304 = idxPagesOH_30 & pageHit;
  assign idxPagesOH_30 = T305[3'h5:1'h0];
  assign T305 = 1'h1 << T306;
  assign T306 = idxPages[6'h1e];
  assign T307 = {T387, T308};
  assign T308 = {T348, T309};
  assign T309 = {T329, T310};
  assign T310 = {T320, T311};
  assign T311 = {T316, T312};
  assign T312 = T313 != 6'h0;
  assign T313 = idxPagesOH_31 & pageHit;
  assign idxPagesOH_31 = T314[3'h5:1'h0];
  assign T314 = 1'h1 << T315;
  assign T315 = idxPages[6'h1f];
  assign T316 = T317 != 6'h0;
  assign T317 = idxPagesOH_32 & pageHit;
  assign idxPagesOH_32 = T318[3'h5:1'h0];
  assign T318 = 1'h1 << T319;
  assign T319 = idxPages[6'h20];
  assign T320 = {T325, T321};
  assign T321 = T322 != 6'h0;
  assign T322 = idxPagesOH_33 & pageHit;
  assign idxPagesOH_33 = T323[3'h5:1'h0];
  assign T323 = 1'h1 << T324;
  assign T324 = idxPages[6'h21];
  assign T325 = T326 != 6'h0;
  assign T326 = idxPagesOH_34 & pageHit;
  assign idxPagesOH_34 = T327[3'h5:1'h0];
  assign T327 = 1'h1 << T328;
  assign T328 = idxPages[6'h22];
  assign T329 = {T339, T330};
  assign T330 = {T335, T331};
  assign T331 = T332 != 6'h0;
  assign T332 = idxPagesOH_35 & pageHit;
  assign idxPagesOH_35 = T333[3'h5:1'h0];
  assign T333 = 1'h1 << T334;
  assign T334 = idxPages[6'h23];
  assign T335 = T336 != 6'h0;
  assign T336 = idxPagesOH_36 & pageHit;
  assign idxPagesOH_36 = T337[3'h5:1'h0];
  assign T337 = 1'h1 << T338;
  assign T338 = idxPages[6'h24];
  assign T339 = {T344, T340};
  assign T340 = T341 != 6'h0;
  assign T341 = idxPagesOH_37 & pageHit;
  assign idxPagesOH_37 = T342[3'h5:1'h0];
  assign T342 = 1'h1 << T343;
  assign T343 = idxPages[6'h25];
  assign T344 = T345 != 6'h0;
  assign T345 = idxPagesOH_38 & pageHit;
  assign idxPagesOH_38 = T346[3'h5:1'h0];
  assign T346 = 1'h1 << T347;
  assign T347 = idxPages[6'h26];
  assign T348 = {T368, T349};
  assign T349 = {T359, T350};
  assign T350 = {T355, T351};
  assign T351 = T352 != 6'h0;
  assign T352 = idxPagesOH_39 & pageHit;
  assign idxPagesOH_39 = T353[3'h5:1'h0];
  assign T353 = 1'h1 << T354;
  assign T354 = idxPages[6'h27];
  assign T355 = T356 != 6'h0;
  assign T356 = idxPagesOH_40 & pageHit;
  assign idxPagesOH_40 = T357[3'h5:1'h0];
  assign T357 = 1'h1 << T358;
  assign T358 = idxPages[6'h28];
  assign T359 = {T364, T360};
  assign T360 = T361 != 6'h0;
  assign T361 = idxPagesOH_41 & pageHit;
  assign idxPagesOH_41 = T362[3'h5:1'h0];
  assign T362 = 1'h1 << T363;
  assign T363 = idxPages[6'h29];
  assign T364 = T365 != 6'h0;
  assign T365 = idxPagesOH_42 & pageHit;
  assign idxPagesOH_42 = T366[3'h5:1'h0];
  assign T366 = 1'h1 << T367;
  assign T367 = idxPages[6'h2a];
  assign T368 = {T378, T369};
  assign T369 = {T374, T370};
  assign T370 = T371 != 6'h0;
  assign T371 = idxPagesOH_43 & pageHit;
  assign idxPagesOH_43 = T372[3'h5:1'h0];
  assign T372 = 1'h1 << T373;
  assign T373 = idxPages[6'h2b];
  assign T374 = T375 != 6'h0;
  assign T375 = idxPagesOH_44 & pageHit;
  assign idxPagesOH_44 = T376[3'h5:1'h0];
  assign T376 = 1'h1 << T377;
  assign T377 = idxPages[6'h2c];
  assign T378 = {T383, T379};
  assign T379 = T380 != 6'h0;
  assign T380 = idxPagesOH_45 & pageHit;
  assign idxPagesOH_45 = T381[3'h5:1'h0];
  assign T381 = 1'h1 << T382;
  assign T382 = idxPages[6'h2d];
  assign T383 = T384 != 6'h0;
  assign T384 = idxPagesOH_46 & pageHit;
  assign idxPagesOH_46 = T385[3'h5:1'h0];
  assign T385 = 1'h1 << T386;
  assign T386 = idxPages[6'h2e];
  assign T387 = {T427, T388};
  assign T388 = {T408, T389};
  assign T389 = {T399, T390};
  assign T390 = {T395, T391};
  assign T391 = T392 != 6'h0;
  assign T392 = idxPagesOH_47 & pageHit;
  assign idxPagesOH_47 = T393[3'h5:1'h0];
  assign T393 = 1'h1 << T394;
  assign T394 = idxPages[6'h2f];
  assign T395 = T396 != 6'h0;
  assign T396 = idxPagesOH_48 & pageHit;
  assign idxPagesOH_48 = T397[3'h5:1'h0];
  assign T397 = 1'h1 << T398;
  assign T398 = idxPages[6'h30];
  assign T399 = {T404, T400};
  assign T400 = T401 != 6'h0;
  assign T401 = idxPagesOH_49 & pageHit;
  assign idxPagesOH_49 = T402[3'h5:1'h0];
  assign T402 = 1'h1 << T403;
  assign T403 = idxPages[6'h31];
  assign T404 = T405 != 6'h0;
  assign T405 = idxPagesOH_50 & pageHit;
  assign idxPagesOH_50 = T406[3'h5:1'h0];
  assign T406 = 1'h1 << T407;
  assign T407 = idxPages[6'h32];
  assign T408 = {T418, T409};
  assign T409 = {T414, T410};
  assign T410 = T411 != 6'h0;
  assign T411 = idxPagesOH_51 & pageHit;
  assign idxPagesOH_51 = T412[3'h5:1'h0];
  assign T412 = 1'h1 << T413;
  assign T413 = idxPages[6'h33];
  assign T414 = T415 != 6'h0;
  assign T415 = idxPagesOH_52 & pageHit;
  assign idxPagesOH_52 = T416[3'h5:1'h0];
  assign T416 = 1'h1 << T417;
  assign T417 = idxPages[6'h34];
  assign T418 = {T423, T419};
  assign T419 = T420 != 6'h0;
  assign T420 = idxPagesOH_53 & pageHit;
  assign idxPagesOH_53 = T421[3'h5:1'h0];
  assign T421 = 1'h1 << T422;
  assign T422 = idxPages[6'h35];
  assign T423 = T424 != 6'h0;
  assign T424 = idxPagesOH_54 & pageHit;
  assign idxPagesOH_54 = T425[3'h5:1'h0];
  assign T425 = 1'h1 << T426;
  assign T426 = idxPages[6'h36];
  assign T427 = {T447, T428};
  assign T428 = {T438, T429};
  assign T429 = {T434, T430};
  assign T430 = T431 != 6'h0;
  assign T431 = idxPagesOH_55 & pageHit;
  assign idxPagesOH_55 = T432[3'h5:1'h0];
  assign T432 = 1'h1 << T433;
  assign T433 = idxPages[6'h37];
  assign T434 = T435 != 6'h0;
  assign T435 = idxPagesOH_56 & pageHit;
  assign idxPagesOH_56 = T436[3'h5:1'h0];
  assign T436 = 1'h1 << T437;
  assign T437 = idxPages[6'h38];
  assign T438 = {T443, T439};
  assign T439 = T440 != 6'h0;
  assign T440 = idxPagesOH_57 & pageHit;
  assign idxPagesOH_57 = T441[3'h5:1'h0];
  assign T441 = 1'h1 << T442;
  assign T442 = idxPages[6'h39];
  assign T443 = T444 != 6'h0;
  assign T444 = idxPagesOH_58 & pageHit;
  assign idxPagesOH_58 = T445[3'h5:1'h0];
  assign T445 = 1'h1 << T446;
  assign T446 = idxPages[6'h3a];
  assign T447 = {T457, T448};
  assign T448 = {T453, T449};
  assign T449 = T450 != 6'h0;
  assign T450 = idxPagesOH_59 & pageHit;
  assign idxPagesOH_59 = T451[3'h5:1'h0];
  assign T451 = 1'h1 << T452;
  assign T452 = idxPages[6'h3b];
  assign T453 = T454 != 6'h0;
  assign T454 = idxPagesOH_60 & pageHit;
  assign idxPagesOH_60 = T455[3'h5:1'h0];
  assign T455 = 1'h1 << T456;
  assign T456 = idxPages[6'h3c];
  assign T457 = T458 != 6'h0;
  assign T458 = idxPagesOH_61 & pageHit;
  assign idxPagesOH_61 = T459[3'h5:1'h0];
  assign T459 = 1'h1 << T460;
  assign T460 = idxPages[6'h3d];
  assign T461 = idxValid & T462;
  assign T462 = T463;
  assign T463 = {T560, T464};
  assign T464 = {T516, T465};
  assign T465 = {T493, T466};
  assign T466 = {T482, T467};
  assign T467 = {T477, T468};
  assign T468 = {T475, T469};
  assign T469 = T471 == T470;
  assign T470 = io_req_bits_addr[4'hb:1'h0];
  assign T471 = idxs[6'h0];
  assign T2305 = R82[4'hb:1'h0];
  assign T473 = R7 & T474;
  assign T474 = T42 < 6'h3e;
  assign T475 = T476 == T470;
  assign T476 = idxs[6'h1];
  assign T477 = {T480, T478};
  assign T478 = T479 == T470;
  assign T479 = idxs[6'h2];
  assign T480 = T481 == T470;
  assign T481 = idxs[6'h3];
  assign T482 = {T488, T483};
  assign T483 = {T486, T484};
  assign T484 = T485 == T470;
  assign T485 = idxs[6'h4];
  assign T486 = T487 == T470;
  assign T487 = idxs[6'h5];
  assign T488 = {T491, T489};
  assign T489 = T490 == T470;
  assign T490 = idxs[6'h6];
  assign T491 = T492 == T470;
  assign T492 = idxs[6'h7];
  assign T493 = {T505, T494};
  assign T494 = {T500, T495};
  assign T495 = {T498, T496};
  assign T496 = T497 == T470;
  assign T497 = idxs[6'h8];
  assign T498 = T499 == T470;
  assign T499 = idxs[6'h9];
  assign T500 = {T503, T501};
  assign T501 = T502 == T470;
  assign T502 = idxs[6'ha];
  assign T503 = T504 == T470;
  assign T504 = idxs[6'hb];
  assign T505 = {T511, T506};
  assign T506 = {T509, T507};
  assign T507 = T508 == T470;
  assign T508 = idxs[6'hc];
  assign T509 = T510 == T470;
  assign T510 = idxs[6'hd];
  assign T511 = {T514, T512};
  assign T512 = T513 == T470;
  assign T513 = idxs[6'he];
  assign T514 = T515 == T470;
  assign T515 = idxs[6'hf];
  assign T516 = {T540, T517};
  assign T517 = {T529, T518};
  assign T518 = {T524, T519};
  assign T519 = {T522, T520};
  assign T520 = T521 == T470;
  assign T521 = idxs[6'h10];
  assign T522 = T523 == T470;
  assign T523 = idxs[6'h11];
  assign T524 = {T527, T525};
  assign T525 = T526 == T470;
  assign T526 = idxs[6'h12];
  assign T527 = T528 == T470;
  assign T528 = idxs[6'h13];
  assign T529 = {T535, T530};
  assign T530 = {T533, T531};
  assign T531 = T532 == T470;
  assign T532 = idxs[6'h14];
  assign T533 = T534 == T470;
  assign T534 = idxs[6'h15];
  assign T535 = {T538, T536};
  assign T536 = T537 == T470;
  assign T537 = idxs[6'h16];
  assign T538 = T539 == T470;
  assign T539 = idxs[6'h17];
  assign T540 = {T552, T541};
  assign T541 = {T547, T542};
  assign T542 = {T545, T543};
  assign T543 = T544 == T470;
  assign T544 = idxs[6'h18];
  assign T545 = T546 == T470;
  assign T546 = idxs[6'h19];
  assign T547 = {T550, T548};
  assign T548 = T549 == T470;
  assign T549 = idxs[6'h1a];
  assign T550 = T551 == T470;
  assign T551 = idxs[6'h1b];
  assign T552 = {T558, T553};
  assign T553 = {T556, T554};
  assign T554 = T555 == T470;
  assign T555 = idxs[6'h1c];
  assign T556 = T557 == T470;
  assign T557 = idxs[6'h1d];
  assign T558 = T559 == T470;
  assign T559 = idxs[6'h1e];
  assign T560 = {T608, T561};
  assign T561 = {T585, T562};
  assign T562 = {T574, T563};
  assign T563 = {T569, T564};
  assign T564 = {T567, T565};
  assign T565 = T566 == T470;
  assign T566 = idxs[6'h1f];
  assign T567 = T568 == T470;
  assign T568 = idxs[6'h20];
  assign T569 = {T572, T570};
  assign T570 = T571 == T470;
  assign T571 = idxs[6'h21];
  assign T572 = T573 == T470;
  assign T573 = idxs[6'h22];
  assign T574 = {T580, T575};
  assign T575 = {T578, T576};
  assign T576 = T577 == T470;
  assign T577 = idxs[6'h23];
  assign T578 = T579 == T470;
  assign T579 = idxs[6'h24];
  assign T580 = {T583, T581};
  assign T581 = T582 == T470;
  assign T582 = idxs[6'h25];
  assign T583 = T584 == T470;
  assign T584 = idxs[6'h26];
  assign T585 = {T597, T586};
  assign T586 = {T592, T587};
  assign T587 = {T590, T588};
  assign T588 = T589 == T470;
  assign T589 = idxs[6'h27];
  assign T590 = T591 == T470;
  assign T591 = idxs[6'h28];
  assign T592 = {T595, T593};
  assign T593 = T594 == T470;
  assign T594 = idxs[6'h29];
  assign T595 = T596 == T470;
  assign T596 = idxs[6'h2a];
  assign T597 = {T603, T598};
  assign T598 = {T601, T599};
  assign T599 = T600 == T470;
  assign T600 = idxs[6'h2b];
  assign T601 = T602 == T470;
  assign T602 = idxs[6'h2c];
  assign T603 = {T606, T604};
  assign T604 = T605 == T470;
  assign T605 = idxs[6'h2d];
  assign T606 = T607 == T470;
  assign T607 = idxs[6'h2e];
  assign T608 = {T632, T609};
  assign T609 = {T621, T610};
  assign T610 = {T616, T611};
  assign T611 = {T614, T612};
  assign T612 = T613 == T470;
  assign T613 = idxs[6'h2f];
  assign T614 = T615 == T470;
  assign T615 = idxs[6'h30];
  assign T616 = {T619, T617};
  assign T617 = T618 == T470;
  assign T618 = idxs[6'h31];
  assign T619 = T620 == T470;
  assign T620 = idxs[6'h32];
  assign T621 = {T627, T622};
  assign T622 = {T625, T623};
  assign T623 = T624 == T470;
  assign T624 = idxs[6'h33];
  assign T625 = T626 == T470;
  assign T626 = idxs[6'h34];
  assign T627 = {T630, T628};
  assign T628 = T629 == T470;
  assign T629 = idxs[6'h35];
  assign T630 = T631 == T470;
  assign T631 = idxs[6'h36];
  assign T632 = {T644, T633};
  assign T633 = {T639, T634};
  assign T634 = {T637, T635};
  assign T635 = T636 == T470;
  assign T636 = idxs[6'h37];
  assign T637 = T638 == T470;
  assign T638 = idxs[6'h38];
  assign T639 = {T642, T640};
  assign T640 = T641 == T470;
  assign T641 = idxs[6'h39];
  assign T642 = T643 == T470;
  assign T643 = idxs[6'h3a];
  assign T644 = {T650, T645};
  assign T645 = {T648, T646};
  assign T646 = T647 == T470;
  assign T647 = idxs[6'h3b];
  assign T648 = T649 == T470;
  assign T649 = idxs[6'h3c];
  assign T650 = T651 == T470;
  assign T651 = idxs[6'h3d];
  assign T2306 = T2307[6'h3d:1'h0];
  assign T2307 = reset ? 64'h0 : T652;
  assign T652 = io_invalidate ? 64'h0 : T653;
  assign T653 = R7 ? T654 : T2308;
  assign T2308 = {2'h0, idxValid};
  assign T654 = T2309 | T655;
  assign T655 = 1'h1 << T42;
  assign T2309 = {2'h0, T656};
  assign T656 = idxValid & T657;
  assign T657 = ~ T658;
  assign T658 = T659;
  assign T659 = {T849, T660};
  assign T660 = {T760, T661};
  assign T661 = {T713, T662};
  assign T662 = {T690, T663};
  assign T663 = {T679, T664};
  assign T664 = {T674, T665};
  assign T665 = T666 != 6'h0;
  assign T666 = pageReplEn & T667;
  assign T667 = idxPagesOH_0 | tgtPagesOH_0;
  assign tgtPagesOH_0 = T668[3'h5:1'h0];
  assign T668 = 1'h1 << T669;
  assign T669 = tgtPages[6'h0];
  assign T2310 = {T2320, T2311};
  assign T2311 = {T2319, T2312};
  assign T2312 = T2313[1'h1:1'h1];
  assign T2313 = T2318 | T2314;
  assign T2314 = T2315[1'h1:1'h0];
  assign T2315 = T2317 | T2316;
  assign T2316 = T671[2'h3:1'h0];
  assign T671 = usePageHit ? pageHit : tgtPageRepl;
  assign T2317 = T671[3'h5:3'h4];
  assign T2318 = T2315[2'h3:2'h2];
  assign T2319 = T2318 != 2'h0;
  assign T2320 = T2317 != 2'h0;
  assign T672 = R7 & T673;
  assign T673 = T42 < 6'h3e;
  assign T674 = T675 != 6'h0;
  assign T675 = pageReplEn & T676;
  assign T676 = idxPagesOH_1 | tgtPagesOH_1;
  assign tgtPagesOH_1 = T677[3'h5:1'h0];
  assign T677 = 1'h1 << T678;
  assign T678 = tgtPages[6'h1];
  assign T679 = {T685, T680};
  assign T680 = T681 != 6'h0;
  assign T681 = pageReplEn & T682;
  assign T682 = idxPagesOH_2 | tgtPagesOH_2;
  assign tgtPagesOH_2 = T683[3'h5:1'h0];
  assign T683 = 1'h1 << T684;
  assign T684 = tgtPages[6'h2];
  assign T685 = T686 != 6'h0;
  assign T686 = pageReplEn & T687;
  assign T687 = idxPagesOH_3 | tgtPagesOH_3;
  assign tgtPagesOH_3 = T688[3'h5:1'h0];
  assign T688 = 1'h1 << T689;
  assign T689 = tgtPages[6'h3];
  assign T690 = {T702, T691};
  assign T691 = {T697, T692};
  assign T692 = T693 != 6'h0;
  assign T693 = pageReplEn & T694;
  assign T694 = idxPagesOH_4 | tgtPagesOH_4;
  assign tgtPagesOH_4 = T695[3'h5:1'h0];
  assign T695 = 1'h1 << T696;
  assign T696 = tgtPages[6'h4];
  assign T697 = T698 != 6'h0;
  assign T698 = pageReplEn & T699;
  assign T699 = idxPagesOH_5 | tgtPagesOH_5;
  assign tgtPagesOH_5 = T700[3'h5:1'h0];
  assign T700 = 1'h1 << T701;
  assign T701 = tgtPages[6'h5];
  assign T702 = {T708, T703};
  assign T703 = T704 != 6'h0;
  assign T704 = pageReplEn & T705;
  assign T705 = idxPagesOH_6 | tgtPagesOH_6;
  assign tgtPagesOH_6 = T706[3'h5:1'h0];
  assign T706 = 1'h1 << T707;
  assign T707 = tgtPages[6'h6];
  assign T708 = T709 != 6'h0;
  assign T709 = pageReplEn & T710;
  assign T710 = idxPagesOH_7 | tgtPagesOH_7;
  assign tgtPagesOH_7 = T711[3'h5:1'h0];
  assign T711 = 1'h1 << T712;
  assign T712 = tgtPages[6'h7];
  assign T713 = {T737, T714};
  assign T714 = {T726, T715};
  assign T715 = {T721, T716};
  assign T716 = T717 != 6'h0;
  assign T717 = pageReplEn & T718;
  assign T718 = idxPagesOH_8 | tgtPagesOH_8;
  assign tgtPagesOH_8 = T719[3'h5:1'h0];
  assign T719 = 1'h1 << T720;
  assign T720 = tgtPages[6'h8];
  assign T721 = T722 != 6'h0;
  assign T722 = pageReplEn & T723;
  assign T723 = idxPagesOH_9 | tgtPagesOH_9;
  assign tgtPagesOH_9 = T724[3'h5:1'h0];
  assign T724 = 1'h1 << T725;
  assign T725 = tgtPages[6'h9];
  assign T726 = {T732, T727};
  assign T727 = T728 != 6'h0;
  assign T728 = pageReplEn & T729;
  assign T729 = idxPagesOH_10 | tgtPagesOH_10;
  assign tgtPagesOH_10 = T730[3'h5:1'h0];
  assign T730 = 1'h1 << T731;
  assign T731 = tgtPages[6'ha];
  assign T732 = T733 != 6'h0;
  assign T733 = pageReplEn & T734;
  assign T734 = idxPagesOH_11 | tgtPagesOH_11;
  assign tgtPagesOH_11 = T735[3'h5:1'h0];
  assign T735 = 1'h1 << T736;
  assign T736 = tgtPages[6'hb];
  assign T737 = {T749, T738};
  assign T738 = {T744, T739};
  assign T739 = T740 != 6'h0;
  assign T740 = pageReplEn & T741;
  assign T741 = idxPagesOH_12 | tgtPagesOH_12;
  assign tgtPagesOH_12 = T742[3'h5:1'h0];
  assign T742 = 1'h1 << T743;
  assign T743 = tgtPages[6'hc];
  assign T744 = T745 != 6'h0;
  assign T745 = pageReplEn & T746;
  assign T746 = idxPagesOH_13 | tgtPagesOH_13;
  assign tgtPagesOH_13 = T747[3'h5:1'h0];
  assign T747 = 1'h1 << T748;
  assign T748 = tgtPages[6'hd];
  assign T749 = {T755, T750};
  assign T750 = T751 != 6'h0;
  assign T751 = pageReplEn & T752;
  assign T752 = idxPagesOH_14 | tgtPagesOH_14;
  assign tgtPagesOH_14 = T753[3'h5:1'h0];
  assign T753 = 1'h1 << T754;
  assign T754 = tgtPages[6'he];
  assign T755 = T756 != 6'h0;
  assign T756 = pageReplEn & T757;
  assign T757 = idxPagesOH_15 | tgtPagesOH_15;
  assign tgtPagesOH_15 = T758[3'h5:1'h0];
  assign T758 = 1'h1 << T759;
  assign T759 = tgtPages[6'hf];
  assign T760 = {T808, T761};
  assign T761 = {T785, T762};
  assign T762 = {T774, T763};
  assign T763 = {T769, T764};
  assign T764 = T765 != 6'h0;
  assign T765 = pageReplEn & T766;
  assign T766 = idxPagesOH_16 | tgtPagesOH_16;
  assign tgtPagesOH_16 = T767[3'h5:1'h0];
  assign T767 = 1'h1 << T768;
  assign T768 = tgtPages[6'h10];
  assign T769 = T770 != 6'h0;
  assign T770 = pageReplEn & T771;
  assign T771 = idxPagesOH_17 | tgtPagesOH_17;
  assign tgtPagesOH_17 = T772[3'h5:1'h0];
  assign T772 = 1'h1 << T773;
  assign T773 = tgtPages[6'h11];
  assign T774 = {T780, T775};
  assign T775 = T776 != 6'h0;
  assign T776 = pageReplEn & T777;
  assign T777 = idxPagesOH_18 | tgtPagesOH_18;
  assign tgtPagesOH_18 = T778[3'h5:1'h0];
  assign T778 = 1'h1 << T779;
  assign T779 = tgtPages[6'h12];
  assign T780 = T781 != 6'h0;
  assign T781 = pageReplEn & T782;
  assign T782 = idxPagesOH_19 | tgtPagesOH_19;
  assign tgtPagesOH_19 = T783[3'h5:1'h0];
  assign T783 = 1'h1 << T784;
  assign T784 = tgtPages[6'h13];
  assign T785 = {T797, T786};
  assign T786 = {T792, T787};
  assign T787 = T788 != 6'h0;
  assign T788 = pageReplEn & T789;
  assign T789 = idxPagesOH_20 | tgtPagesOH_20;
  assign tgtPagesOH_20 = T790[3'h5:1'h0];
  assign T790 = 1'h1 << T791;
  assign T791 = tgtPages[6'h14];
  assign T792 = T793 != 6'h0;
  assign T793 = pageReplEn & T794;
  assign T794 = idxPagesOH_21 | tgtPagesOH_21;
  assign tgtPagesOH_21 = T795[3'h5:1'h0];
  assign T795 = 1'h1 << T796;
  assign T796 = tgtPages[6'h15];
  assign T797 = {T803, T798};
  assign T798 = T799 != 6'h0;
  assign T799 = pageReplEn & T800;
  assign T800 = idxPagesOH_22 | tgtPagesOH_22;
  assign tgtPagesOH_22 = T801[3'h5:1'h0];
  assign T801 = 1'h1 << T802;
  assign T802 = tgtPages[6'h16];
  assign T803 = T804 != 6'h0;
  assign T804 = pageReplEn & T805;
  assign T805 = idxPagesOH_23 | tgtPagesOH_23;
  assign tgtPagesOH_23 = T806[3'h5:1'h0];
  assign T806 = 1'h1 << T807;
  assign T807 = tgtPages[6'h17];
  assign T808 = {T832, T809};
  assign T809 = {T821, T810};
  assign T810 = {T816, T811};
  assign T811 = T812 != 6'h0;
  assign T812 = pageReplEn & T813;
  assign T813 = idxPagesOH_24 | tgtPagesOH_24;
  assign tgtPagesOH_24 = T814[3'h5:1'h0];
  assign T814 = 1'h1 << T815;
  assign T815 = tgtPages[6'h18];
  assign T816 = T817 != 6'h0;
  assign T817 = pageReplEn & T818;
  assign T818 = idxPagesOH_25 | tgtPagesOH_25;
  assign tgtPagesOH_25 = T819[3'h5:1'h0];
  assign T819 = 1'h1 << T820;
  assign T820 = tgtPages[6'h19];
  assign T821 = {T827, T822};
  assign T822 = T823 != 6'h0;
  assign T823 = pageReplEn & T824;
  assign T824 = idxPagesOH_26 | tgtPagesOH_26;
  assign tgtPagesOH_26 = T825[3'h5:1'h0];
  assign T825 = 1'h1 << T826;
  assign T826 = tgtPages[6'h1a];
  assign T827 = T828 != 6'h0;
  assign T828 = pageReplEn & T829;
  assign T829 = idxPagesOH_27 | tgtPagesOH_27;
  assign tgtPagesOH_27 = T830[3'h5:1'h0];
  assign T830 = 1'h1 << T831;
  assign T831 = tgtPages[6'h1b];
  assign T832 = {T844, T833};
  assign T833 = {T839, T834};
  assign T834 = T835 != 6'h0;
  assign T835 = pageReplEn & T836;
  assign T836 = idxPagesOH_28 | tgtPagesOH_28;
  assign tgtPagesOH_28 = T837[3'h5:1'h0];
  assign T837 = 1'h1 << T838;
  assign T838 = tgtPages[6'h1c];
  assign T839 = T840 != 6'h0;
  assign T840 = pageReplEn & T841;
  assign T841 = idxPagesOH_29 | tgtPagesOH_29;
  assign tgtPagesOH_29 = T842[3'h5:1'h0];
  assign T842 = 1'h1 << T843;
  assign T843 = tgtPages[6'h1d];
  assign T844 = T845 != 6'h0;
  assign T845 = pageReplEn & T846;
  assign T846 = idxPagesOH_30 | tgtPagesOH_30;
  assign tgtPagesOH_30 = T847[3'h5:1'h0];
  assign T847 = 1'h1 << T848;
  assign T848 = tgtPages[6'h1e];
  assign T849 = {T945, T850};
  assign T850 = {T898, T851};
  assign T851 = {T875, T852};
  assign T852 = {T864, T853};
  assign T853 = {T859, T854};
  assign T854 = T855 != 6'h0;
  assign T855 = pageReplEn & T856;
  assign T856 = idxPagesOH_31 | tgtPagesOH_31;
  assign tgtPagesOH_31 = T857[3'h5:1'h0];
  assign T857 = 1'h1 << T858;
  assign T858 = tgtPages[6'h1f];
  assign T859 = T860 != 6'h0;
  assign T860 = pageReplEn & T861;
  assign T861 = idxPagesOH_32 | tgtPagesOH_32;
  assign tgtPagesOH_32 = T862[3'h5:1'h0];
  assign T862 = 1'h1 << T863;
  assign T863 = tgtPages[6'h20];
  assign T864 = {T870, T865};
  assign T865 = T866 != 6'h0;
  assign T866 = pageReplEn & T867;
  assign T867 = idxPagesOH_33 | tgtPagesOH_33;
  assign tgtPagesOH_33 = T868[3'h5:1'h0];
  assign T868 = 1'h1 << T869;
  assign T869 = tgtPages[6'h21];
  assign T870 = T871 != 6'h0;
  assign T871 = pageReplEn & T872;
  assign T872 = idxPagesOH_34 | tgtPagesOH_34;
  assign tgtPagesOH_34 = T873[3'h5:1'h0];
  assign T873 = 1'h1 << T874;
  assign T874 = tgtPages[6'h22];
  assign T875 = {T887, T876};
  assign T876 = {T882, T877};
  assign T877 = T878 != 6'h0;
  assign T878 = pageReplEn & T879;
  assign T879 = idxPagesOH_35 | tgtPagesOH_35;
  assign tgtPagesOH_35 = T880[3'h5:1'h0];
  assign T880 = 1'h1 << T881;
  assign T881 = tgtPages[6'h23];
  assign T882 = T883 != 6'h0;
  assign T883 = pageReplEn & T884;
  assign T884 = idxPagesOH_36 | tgtPagesOH_36;
  assign tgtPagesOH_36 = T885[3'h5:1'h0];
  assign T885 = 1'h1 << T886;
  assign T886 = tgtPages[6'h24];
  assign T887 = {T893, T888};
  assign T888 = T889 != 6'h0;
  assign T889 = pageReplEn & T890;
  assign T890 = idxPagesOH_37 | tgtPagesOH_37;
  assign tgtPagesOH_37 = T891[3'h5:1'h0];
  assign T891 = 1'h1 << T892;
  assign T892 = tgtPages[6'h25];
  assign T893 = T894 != 6'h0;
  assign T894 = pageReplEn & T895;
  assign T895 = idxPagesOH_38 | tgtPagesOH_38;
  assign tgtPagesOH_38 = T896[3'h5:1'h0];
  assign T896 = 1'h1 << T897;
  assign T897 = tgtPages[6'h26];
  assign T898 = {T922, T899};
  assign T899 = {T911, T900};
  assign T900 = {T906, T901};
  assign T901 = T902 != 6'h0;
  assign T902 = pageReplEn & T903;
  assign T903 = idxPagesOH_39 | tgtPagesOH_39;
  assign tgtPagesOH_39 = T904[3'h5:1'h0];
  assign T904 = 1'h1 << T905;
  assign T905 = tgtPages[6'h27];
  assign T906 = T907 != 6'h0;
  assign T907 = pageReplEn & T908;
  assign T908 = idxPagesOH_40 | tgtPagesOH_40;
  assign tgtPagesOH_40 = T909[3'h5:1'h0];
  assign T909 = 1'h1 << T910;
  assign T910 = tgtPages[6'h28];
  assign T911 = {T917, T912};
  assign T912 = T913 != 6'h0;
  assign T913 = pageReplEn & T914;
  assign T914 = idxPagesOH_41 | tgtPagesOH_41;
  assign tgtPagesOH_41 = T915[3'h5:1'h0];
  assign T915 = 1'h1 << T916;
  assign T916 = tgtPages[6'h29];
  assign T917 = T918 != 6'h0;
  assign T918 = pageReplEn & T919;
  assign T919 = idxPagesOH_42 | tgtPagesOH_42;
  assign tgtPagesOH_42 = T920[3'h5:1'h0];
  assign T920 = 1'h1 << T921;
  assign T921 = tgtPages[6'h2a];
  assign T922 = {T934, T923};
  assign T923 = {T929, T924};
  assign T924 = T925 != 6'h0;
  assign T925 = pageReplEn & T926;
  assign T926 = idxPagesOH_43 | tgtPagesOH_43;
  assign tgtPagesOH_43 = T927[3'h5:1'h0];
  assign T927 = 1'h1 << T928;
  assign T928 = tgtPages[6'h2b];
  assign T929 = T930 != 6'h0;
  assign T930 = pageReplEn & T931;
  assign T931 = idxPagesOH_44 | tgtPagesOH_44;
  assign tgtPagesOH_44 = T932[3'h5:1'h0];
  assign T932 = 1'h1 << T933;
  assign T933 = tgtPages[6'h2c];
  assign T934 = {T940, T935};
  assign T935 = T936 != 6'h0;
  assign T936 = pageReplEn & T937;
  assign T937 = idxPagesOH_45 | tgtPagesOH_45;
  assign tgtPagesOH_45 = T938[3'h5:1'h0];
  assign T938 = 1'h1 << T939;
  assign T939 = tgtPages[6'h2d];
  assign T940 = T941 != 6'h0;
  assign T941 = pageReplEn & T942;
  assign T942 = idxPagesOH_46 | tgtPagesOH_46;
  assign tgtPagesOH_46 = T943[3'h5:1'h0];
  assign T943 = 1'h1 << T944;
  assign T944 = tgtPages[6'h2e];
  assign T945 = {T993, T946};
  assign T946 = {T970, T947};
  assign T947 = {T959, T948};
  assign T948 = {T954, T949};
  assign T949 = T950 != 6'h0;
  assign T950 = pageReplEn & T951;
  assign T951 = idxPagesOH_47 | tgtPagesOH_47;
  assign tgtPagesOH_47 = T952[3'h5:1'h0];
  assign T952 = 1'h1 << T953;
  assign T953 = tgtPages[6'h2f];
  assign T954 = T955 != 6'h0;
  assign T955 = pageReplEn & T956;
  assign T956 = idxPagesOH_48 | tgtPagesOH_48;
  assign tgtPagesOH_48 = T957[3'h5:1'h0];
  assign T957 = 1'h1 << T958;
  assign T958 = tgtPages[6'h30];
  assign T959 = {T965, T960};
  assign T960 = T961 != 6'h0;
  assign T961 = pageReplEn & T962;
  assign T962 = idxPagesOH_49 | tgtPagesOH_49;
  assign tgtPagesOH_49 = T963[3'h5:1'h0];
  assign T963 = 1'h1 << T964;
  assign T964 = tgtPages[6'h31];
  assign T965 = T966 != 6'h0;
  assign T966 = pageReplEn & T967;
  assign T967 = idxPagesOH_50 | tgtPagesOH_50;
  assign tgtPagesOH_50 = T968[3'h5:1'h0];
  assign T968 = 1'h1 << T969;
  assign T969 = tgtPages[6'h32];
  assign T970 = {T982, T971};
  assign T971 = {T977, T972};
  assign T972 = T973 != 6'h0;
  assign T973 = pageReplEn & T974;
  assign T974 = idxPagesOH_51 | tgtPagesOH_51;
  assign tgtPagesOH_51 = T975[3'h5:1'h0];
  assign T975 = 1'h1 << T976;
  assign T976 = tgtPages[6'h33];
  assign T977 = T978 != 6'h0;
  assign T978 = pageReplEn & T979;
  assign T979 = idxPagesOH_52 | tgtPagesOH_52;
  assign tgtPagesOH_52 = T980[3'h5:1'h0];
  assign T980 = 1'h1 << T981;
  assign T981 = tgtPages[6'h34];
  assign T982 = {T988, T983};
  assign T983 = T984 != 6'h0;
  assign T984 = pageReplEn & T985;
  assign T985 = idxPagesOH_53 | tgtPagesOH_53;
  assign tgtPagesOH_53 = T986[3'h5:1'h0];
  assign T986 = 1'h1 << T987;
  assign T987 = tgtPages[6'h35];
  assign T988 = T989 != 6'h0;
  assign T989 = pageReplEn & T990;
  assign T990 = idxPagesOH_54 | tgtPagesOH_54;
  assign tgtPagesOH_54 = T991[3'h5:1'h0];
  assign T991 = 1'h1 << T992;
  assign T992 = tgtPages[6'h36];
  assign T993 = {T1017, T994};
  assign T994 = {T1006, T995};
  assign T995 = {T1001, T996};
  assign T996 = T997 != 6'h0;
  assign T997 = pageReplEn & T998;
  assign T998 = idxPagesOH_55 | tgtPagesOH_55;
  assign tgtPagesOH_55 = T999[3'h5:1'h0];
  assign T999 = 1'h1 << T1000;
  assign T1000 = tgtPages[6'h37];
  assign T1001 = T1002 != 6'h0;
  assign T1002 = pageReplEn & T1003;
  assign T1003 = idxPagesOH_56 | tgtPagesOH_56;
  assign tgtPagesOH_56 = T1004[3'h5:1'h0];
  assign T1004 = 1'h1 << T1005;
  assign T1005 = tgtPages[6'h38];
  assign T1006 = {T1012, T1007};
  assign T1007 = T1008 != 6'h0;
  assign T1008 = pageReplEn & T1009;
  assign T1009 = idxPagesOH_57 | tgtPagesOH_57;
  assign tgtPagesOH_57 = T1010[3'h5:1'h0];
  assign T1010 = 1'h1 << T1011;
  assign T1011 = tgtPages[6'h39];
  assign T1012 = T1013 != 6'h0;
  assign T1013 = pageReplEn & T1014;
  assign T1014 = idxPagesOH_58 | tgtPagesOH_58;
  assign tgtPagesOH_58 = T1015[3'h5:1'h0];
  assign T1015 = 1'h1 << T1016;
  assign T1016 = tgtPages[6'h3a];
  assign T1017 = {T1029, T1018};
  assign T1018 = {T1024, T1019};
  assign T1019 = T1020 != 6'h0;
  assign T1020 = pageReplEn & T1021;
  assign T1021 = idxPagesOH_59 | tgtPagesOH_59;
  assign tgtPagesOH_59 = T1022[3'h5:1'h0];
  assign T1022 = 1'h1 << T1023;
  assign T1023 = tgtPages[6'h3b];
  assign T1024 = T1025 != 6'h0;
  assign T1025 = pageReplEn & T1026;
  assign T1026 = idxPagesOH_60 | tgtPagesOH_60;
  assign tgtPagesOH_60 = T1027[3'h5:1'h0];
  assign T1027 = 1'h1 << T1028;
  assign T1028 = tgtPages[6'h3c];
  assign T1029 = T1030 != 6'h0;
  assign T1030 = pageReplEn & T1031;
  assign T1031 = idxPagesOH_61 | tgtPagesOH_61;
  assign tgtPagesOH_61 = T1032[3'h5:1'h0];
  assign T1032 = 1'h1 << T1033;
  assign T1033 = tgtPages[6'h3d];
  assign T1034 = T1040 | T1035;
  assign T1035 = T1039 ? isJump_60 : 1'h0;
  assign T1036 = T1037 ? R36 : isJump_60;
  assign T1037 = R7 & T1038;
  assign T1038 = T40[6'h3c:6'h3c];
  assign T1039 = hits[6'h3c:6'h3c];
  assign T1040 = T1046 | T1041;
  assign T1041 = T1045 ? isJump_59 : 1'h0;
  assign T1042 = T1043 ? R36 : isJump_59;
  assign T1043 = R7 & T1044;
  assign T1044 = T40[6'h3b:6'h3b];
  assign T1045 = hits[6'h3b:6'h3b];
  assign T1046 = T1052 | T1047;
  assign T1047 = T1051 ? isJump_58 : 1'h0;
  assign T1048 = T1049 ? R36 : isJump_58;
  assign T1049 = R7 & T1050;
  assign T1050 = T40[6'h3a:6'h3a];
  assign T1051 = hits[6'h3a:6'h3a];
  assign T1052 = T1058 | T1053;
  assign T1053 = T1057 ? isJump_57 : 1'h0;
  assign T1054 = T1055 ? R36 : isJump_57;
  assign T1055 = R7 & T1056;
  assign T1056 = T40[6'h39:6'h39];
  assign T1057 = hits[6'h39:6'h39];
  assign T1058 = T1064 | T1059;
  assign T1059 = T1063 ? isJump_56 : 1'h0;
  assign T1060 = T1061 ? R36 : isJump_56;
  assign T1061 = R7 & T1062;
  assign T1062 = T40[6'h38:6'h38];
  assign T1063 = hits[6'h38:6'h38];
  assign T1064 = T1070 | T1065;
  assign T1065 = T1069 ? isJump_55 : 1'h0;
  assign T1066 = T1067 ? R36 : isJump_55;
  assign T1067 = R7 & T1068;
  assign T1068 = T40[6'h37:6'h37];
  assign T1069 = hits[6'h37:6'h37];
  assign T1070 = T1076 | T1071;
  assign T1071 = T1075 ? isJump_54 : 1'h0;
  assign T1072 = T1073 ? R36 : isJump_54;
  assign T1073 = R7 & T1074;
  assign T1074 = T40[6'h36:6'h36];
  assign T1075 = hits[6'h36:6'h36];
  assign T1076 = T1082 | T1077;
  assign T1077 = T1081 ? isJump_53 : 1'h0;
  assign T1078 = T1079 ? R36 : isJump_53;
  assign T1079 = R7 & T1080;
  assign T1080 = T40[6'h35:6'h35];
  assign T1081 = hits[6'h35:6'h35];
  assign T1082 = T1088 | T1083;
  assign T1083 = T1087 ? isJump_52 : 1'h0;
  assign T1084 = T1085 ? R36 : isJump_52;
  assign T1085 = R7 & T1086;
  assign T1086 = T40[6'h34:6'h34];
  assign T1087 = hits[6'h34:6'h34];
  assign T1088 = T1094 | T1089;
  assign T1089 = T1093 ? isJump_51 : 1'h0;
  assign T1090 = T1091 ? R36 : isJump_51;
  assign T1091 = R7 & T1092;
  assign T1092 = T40[6'h33:6'h33];
  assign T1093 = hits[6'h33:6'h33];
  assign T1094 = T1100 | T1095;
  assign T1095 = T1099 ? isJump_50 : 1'h0;
  assign T1096 = T1097 ? R36 : isJump_50;
  assign T1097 = R7 & T1098;
  assign T1098 = T40[6'h32:6'h32];
  assign T1099 = hits[6'h32:6'h32];
  assign T1100 = T1106 | T1101;
  assign T1101 = T1105 ? isJump_49 : 1'h0;
  assign T1102 = T1103 ? R36 : isJump_49;
  assign T1103 = R7 & T1104;
  assign T1104 = T40[6'h31:6'h31];
  assign T1105 = hits[6'h31:6'h31];
  assign T1106 = T1112 | T1107;
  assign T1107 = T1111 ? isJump_48 : 1'h0;
  assign T1108 = T1109 ? R36 : isJump_48;
  assign T1109 = R7 & T1110;
  assign T1110 = T40[6'h30:6'h30];
  assign T1111 = hits[6'h30:6'h30];
  assign T1112 = T1118 | T1113;
  assign T1113 = T1117 ? isJump_47 : 1'h0;
  assign T1114 = T1115 ? R36 : isJump_47;
  assign T1115 = R7 & T1116;
  assign T1116 = T40[6'h2f:6'h2f];
  assign T1117 = hits[6'h2f:6'h2f];
  assign T1118 = T1124 | T1119;
  assign T1119 = T1123 ? isJump_46 : 1'h0;
  assign T1120 = T1121 ? R36 : isJump_46;
  assign T1121 = R7 & T1122;
  assign T1122 = T40[6'h2e:6'h2e];
  assign T1123 = hits[6'h2e:6'h2e];
  assign T1124 = T1130 | T1125;
  assign T1125 = T1129 ? isJump_45 : 1'h0;
  assign T1126 = T1127 ? R36 : isJump_45;
  assign T1127 = R7 & T1128;
  assign T1128 = T40[6'h2d:6'h2d];
  assign T1129 = hits[6'h2d:6'h2d];
  assign T1130 = T1136 | T1131;
  assign T1131 = T1135 ? isJump_44 : 1'h0;
  assign T1132 = T1133 ? R36 : isJump_44;
  assign T1133 = R7 & T1134;
  assign T1134 = T40[6'h2c:6'h2c];
  assign T1135 = hits[6'h2c:6'h2c];
  assign T1136 = T1142 | T1137;
  assign T1137 = T1141 ? isJump_43 : 1'h0;
  assign T1138 = T1139 ? R36 : isJump_43;
  assign T1139 = R7 & T1140;
  assign T1140 = T40[6'h2b:6'h2b];
  assign T1141 = hits[6'h2b:6'h2b];
  assign T1142 = T1148 | T1143;
  assign T1143 = T1147 ? isJump_42 : 1'h0;
  assign T1144 = T1145 ? R36 : isJump_42;
  assign T1145 = R7 & T1146;
  assign T1146 = T40[6'h2a:6'h2a];
  assign T1147 = hits[6'h2a:6'h2a];
  assign T1148 = T1154 | T1149;
  assign T1149 = T1153 ? isJump_41 : 1'h0;
  assign T1150 = T1151 ? R36 : isJump_41;
  assign T1151 = R7 & T1152;
  assign T1152 = T40[6'h29:6'h29];
  assign T1153 = hits[6'h29:6'h29];
  assign T1154 = T1160 | T1155;
  assign T1155 = T1159 ? isJump_40 : 1'h0;
  assign T1156 = T1157 ? R36 : isJump_40;
  assign T1157 = R7 & T1158;
  assign T1158 = T40[6'h28:6'h28];
  assign T1159 = hits[6'h28:6'h28];
  assign T1160 = T1166 | T1161;
  assign T1161 = T1165 ? isJump_39 : 1'h0;
  assign T1162 = T1163 ? R36 : isJump_39;
  assign T1163 = R7 & T1164;
  assign T1164 = T40[6'h27:6'h27];
  assign T1165 = hits[6'h27:6'h27];
  assign T1166 = T1172 | T1167;
  assign T1167 = T1171 ? isJump_38 : 1'h0;
  assign T1168 = T1169 ? R36 : isJump_38;
  assign T1169 = R7 & T1170;
  assign T1170 = T40[6'h26:6'h26];
  assign T1171 = hits[6'h26:6'h26];
  assign T1172 = T1178 | T1173;
  assign T1173 = T1177 ? isJump_37 : 1'h0;
  assign T1174 = T1175 ? R36 : isJump_37;
  assign T1175 = R7 & T1176;
  assign T1176 = T40[6'h25:6'h25];
  assign T1177 = hits[6'h25:6'h25];
  assign T1178 = T1184 | T1179;
  assign T1179 = T1183 ? isJump_36 : 1'h0;
  assign T1180 = T1181 ? R36 : isJump_36;
  assign T1181 = R7 & T1182;
  assign T1182 = T40[6'h24:6'h24];
  assign T1183 = hits[6'h24:6'h24];
  assign T1184 = T1190 | T1185;
  assign T1185 = T1189 ? isJump_35 : 1'h0;
  assign T1186 = T1187 ? R36 : isJump_35;
  assign T1187 = R7 & T1188;
  assign T1188 = T40[6'h23:6'h23];
  assign T1189 = hits[6'h23:6'h23];
  assign T1190 = T1196 | T1191;
  assign T1191 = T1195 ? isJump_34 : 1'h0;
  assign T1192 = T1193 ? R36 : isJump_34;
  assign T1193 = R7 & T1194;
  assign T1194 = T40[6'h22:6'h22];
  assign T1195 = hits[6'h22:6'h22];
  assign T1196 = T1202 | T1197;
  assign T1197 = T1201 ? isJump_33 : 1'h0;
  assign T1198 = T1199 ? R36 : isJump_33;
  assign T1199 = R7 & T1200;
  assign T1200 = T40[6'h21:6'h21];
  assign T1201 = hits[6'h21:6'h21];
  assign T1202 = T1208 | T1203;
  assign T1203 = T1207 ? isJump_32 : 1'h0;
  assign T1204 = T1205 ? R36 : isJump_32;
  assign T1205 = R7 & T1206;
  assign T1206 = T40[6'h20:6'h20];
  assign T1207 = hits[6'h20:6'h20];
  assign T1208 = T1214 | T1209;
  assign T1209 = T1213 ? isJump_31 : 1'h0;
  assign T1210 = T1211 ? R36 : isJump_31;
  assign T1211 = R7 & T1212;
  assign T1212 = T40[5'h1f:5'h1f];
  assign T1213 = hits[5'h1f:5'h1f];
  assign T1214 = T1220 | T1215;
  assign T1215 = T1219 ? isJump_30 : 1'h0;
  assign T1216 = T1217 ? R36 : isJump_30;
  assign T1217 = R7 & T1218;
  assign T1218 = T40[5'h1e:5'h1e];
  assign T1219 = hits[5'h1e:5'h1e];
  assign T1220 = T1226 | T1221;
  assign T1221 = T1225 ? isJump_29 : 1'h0;
  assign T1222 = T1223 ? R36 : isJump_29;
  assign T1223 = R7 & T1224;
  assign T1224 = T40[5'h1d:5'h1d];
  assign T1225 = hits[5'h1d:5'h1d];
  assign T1226 = T1232 | T1227;
  assign T1227 = T1231 ? isJump_28 : 1'h0;
  assign T1228 = T1229 ? R36 : isJump_28;
  assign T1229 = R7 & T1230;
  assign T1230 = T40[5'h1c:5'h1c];
  assign T1231 = hits[5'h1c:5'h1c];
  assign T1232 = T1238 | T1233;
  assign T1233 = T1237 ? isJump_27 : 1'h0;
  assign T1234 = T1235 ? R36 : isJump_27;
  assign T1235 = R7 & T1236;
  assign T1236 = T40[5'h1b:5'h1b];
  assign T1237 = hits[5'h1b:5'h1b];
  assign T1238 = T1244 | T1239;
  assign T1239 = T1243 ? isJump_26 : 1'h0;
  assign T1240 = T1241 ? R36 : isJump_26;
  assign T1241 = R7 & T1242;
  assign T1242 = T40[5'h1a:5'h1a];
  assign T1243 = hits[5'h1a:5'h1a];
  assign T1244 = T1250 | T1245;
  assign T1245 = T1249 ? isJump_25 : 1'h0;
  assign T1246 = T1247 ? R36 : isJump_25;
  assign T1247 = R7 & T1248;
  assign T1248 = T40[5'h19:5'h19];
  assign T1249 = hits[5'h19:5'h19];
  assign T1250 = T1256 | T1251;
  assign T1251 = T1255 ? isJump_24 : 1'h0;
  assign T1252 = T1253 ? R36 : isJump_24;
  assign T1253 = R7 & T1254;
  assign T1254 = T40[5'h18:5'h18];
  assign T1255 = hits[5'h18:5'h18];
  assign T1256 = T1262 | T1257;
  assign T1257 = T1261 ? isJump_23 : 1'h0;
  assign T1258 = T1259 ? R36 : isJump_23;
  assign T1259 = R7 & T1260;
  assign T1260 = T40[5'h17:5'h17];
  assign T1261 = hits[5'h17:5'h17];
  assign T1262 = T1268 | T1263;
  assign T1263 = T1267 ? isJump_22 : 1'h0;
  assign T1264 = T1265 ? R36 : isJump_22;
  assign T1265 = R7 & T1266;
  assign T1266 = T40[5'h16:5'h16];
  assign T1267 = hits[5'h16:5'h16];
  assign T1268 = T1274 | T1269;
  assign T1269 = T1273 ? isJump_21 : 1'h0;
  assign T1270 = T1271 ? R36 : isJump_21;
  assign T1271 = R7 & T1272;
  assign T1272 = T40[5'h15:5'h15];
  assign T1273 = hits[5'h15:5'h15];
  assign T1274 = T1280 | T1275;
  assign T1275 = T1279 ? isJump_20 : 1'h0;
  assign T1276 = T1277 ? R36 : isJump_20;
  assign T1277 = R7 & T1278;
  assign T1278 = T40[5'h14:5'h14];
  assign T1279 = hits[5'h14:5'h14];
  assign T1280 = T1286 | T1281;
  assign T1281 = T1285 ? isJump_19 : 1'h0;
  assign T1282 = T1283 ? R36 : isJump_19;
  assign T1283 = R7 & T1284;
  assign T1284 = T40[5'h13:5'h13];
  assign T1285 = hits[5'h13:5'h13];
  assign T1286 = T1292 | T1287;
  assign T1287 = T1291 ? isJump_18 : 1'h0;
  assign T1288 = T1289 ? R36 : isJump_18;
  assign T1289 = R7 & T1290;
  assign T1290 = T40[5'h12:5'h12];
  assign T1291 = hits[5'h12:5'h12];
  assign T1292 = T1298 | T1293;
  assign T1293 = T1297 ? isJump_17 : 1'h0;
  assign T1294 = T1295 ? R36 : isJump_17;
  assign T1295 = R7 & T1296;
  assign T1296 = T40[5'h11:5'h11];
  assign T1297 = hits[5'h11:5'h11];
  assign T1298 = T1304 | T1299;
  assign T1299 = T1303 ? isJump_16 : 1'h0;
  assign T1300 = T1301 ? R36 : isJump_16;
  assign T1301 = R7 & T1302;
  assign T1302 = T40[5'h10:5'h10];
  assign T1303 = hits[5'h10:5'h10];
  assign T1304 = T1310 | T1305;
  assign T1305 = T1309 ? isJump_15 : 1'h0;
  assign T1306 = T1307 ? R36 : isJump_15;
  assign T1307 = R7 & T1308;
  assign T1308 = T40[4'hf:4'hf];
  assign T1309 = hits[4'hf:4'hf];
  assign T1310 = T1316 | T1311;
  assign T1311 = T1315 ? isJump_14 : 1'h0;
  assign T1312 = T1313 ? R36 : isJump_14;
  assign T1313 = R7 & T1314;
  assign T1314 = T40[4'he:4'he];
  assign T1315 = hits[4'he:4'he];
  assign T1316 = T1322 | T1317;
  assign T1317 = T1321 ? isJump_13 : 1'h0;
  assign T1318 = T1319 ? R36 : isJump_13;
  assign T1319 = R7 & T1320;
  assign T1320 = T40[4'hd:4'hd];
  assign T1321 = hits[4'hd:4'hd];
  assign T1322 = T1328 | T1323;
  assign T1323 = T1327 ? isJump_12 : 1'h0;
  assign T1324 = T1325 ? R36 : isJump_12;
  assign T1325 = R7 & T1326;
  assign T1326 = T40[4'hc:4'hc];
  assign T1327 = hits[4'hc:4'hc];
  assign T1328 = T1334 | T1329;
  assign T1329 = T1333 ? isJump_11 : 1'h0;
  assign T1330 = T1331 ? R36 : isJump_11;
  assign T1331 = R7 & T1332;
  assign T1332 = T40[4'hb:4'hb];
  assign T1333 = hits[4'hb:4'hb];
  assign T1334 = T1340 | T1335;
  assign T1335 = T1339 ? isJump_10 : 1'h0;
  assign T1336 = T1337 ? R36 : isJump_10;
  assign T1337 = R7 & T1338;
  assign T1338 = T40[4'ha:4'ha];
  assign T1339 = hits[4'ha:4'ha];
  assign T1340 = T1346 | T1341;
  assign T1341 = T1345 ? isJump_9 : 1'h0;
  assign T1342 = T1343 ? R36 : isJump_9;
  assign T1343 = R7 & T1344;
  assign T1344 = T40[4'h9:4'h9];
  assign T1345 = hits[4'h9:4'h9];
  assign T1346 = T1352 | T1347;
  assign T1347 = T1351 ? isJump_8 : 1'h0;
  assign T1348 = T1349 ? R36 : isJump_8;
  assign T1349 = R7 & T1350;
  assign T1350 = T40[4'h8:4'h8];
  assign T1351 = hits[4'h8:4'h8];
  assign T1352 = T1358 | T1353;
  assign T1353 = T1357 ? isJump_7 : 1'h0;
  assign T1354 = T1355 ? R36 : isJump_7;
  assign T1355 = R7 & T1356;
  assign T1356 = T40[3'h7:3'h7];
  assign T1357 = hits[3'h7:3'h7];
  assign T1358 = T1364 | T1359;
  assign T1359 = T1363 ? isJump_6 : 1'h0;
  assign T1360 = T1361 ? R36 : isJump_6;
  assign T1361 = R7 & T1362;
  assign T1362 = T40[3'h6:3'h6];
  assign T1363 = hits[3'h6:3'h6];
  assign T1364 = T1370 | T1365;
  assign T1365 = T1369 ? isJump_5 : 1'h0;
  assign T1366 = T1367 ? R36 : isJump_5;
  assign T1367 = R7 & T1368;
  assign T1368 = T40[3'h5:3'h5];
  assign T1369 = hits[3'h5:3'h5];
  assign T1370 = T1376 | T1371;
  assign T1371 = T1375 ? isJump_4 : 1'h0;
  assign T1372 = T1373 ? R36 : isJump_4;
  assign T1373 = R7 & T1374;
  assign T1374 = T40[3'h4:3'h4];
  assign T1375 = hits[3'h4:3'h4];
  assign T1376 = T1382 | T1377;
  assign T1377 = T1381 ? isJump_3 : 1'h0;
  assign T1378 = T1379 ? R36 : isJump_3;
  assign T1379 = R7 & T1380;
  assign T1380 = T40[2'h3:2'h3];
  assign T1381 = hits[2'h3:2'h3];
  assign T1382 = T1388 | T1383;
  assign T1383 = T1387 ? isJump_2 : 1'h0;
  assign T1384 = T1385 ? R36 : isJump_2;
  assign T1385 = R7 & T1386;
  assign T1386 = T40[2'h2:2'h2];
  assign T1387 = hits[2'h2:2'h2];
  assign T1388 = T1394 | T1389;
  assign T1389 = T1393 ? isJump_1 : 1'h0;
  assign T1390 = T1391 ? R36 : isJump_1;
  assign T1391 = R7 & T1392;
  assign T1392 = T40[1'h1:1'h1];
  assign T1393 = hits[1'h1:1'h1];
  assign T1394 = T1398 ? isJump_0 : 1'h0;
  assign T1395 = T1396 ? R36 : isJump_0;
  assign T1396 = R7 & T1397;
  assign T1397 = T40[1'h0:1'h0];
  assign T1398 = hits[1'h0:1'h0];
  assign T1399 = io_req_valid & io_resp_valid;
  assign T1400 = {io_bht_update_bits_taken, T1401};
  assign T1401 = io_bht_update_bits_prediction_bits_bht_history[3'h6:1'h1];
  assign T1402 = T21 & io_bht_update_bits_mispredict;
  assign T1403 = io_req_bits_addr[4'h8:2'h2];
  assign io_resp_bits_bht_history = T1404;
  assign T1404 = R25;
  assign io_resp_bits_entry = T2321;
  assign T2321 = {T2346, T2322};
  assign T2322 = {T2345, T2323};
  assign T2323 = {T2344, T2324};
  assign T2324 = {T2343, T2325};
  assign T2325 = {T2342, T2326};
  assign T2326 = T2327[1'h1:1'h1];
  assign T2327 = T2341 | T2328;
  assign T2328 = T2329[1'h1:1'h0];
  assign T2329 = T2340 | T2330;
  assign T2330 = T2331[2'h3:1'h0];
  assign T2331 = T2339 | T2332;
  assign T2332 = T2333[3'h7:1'h0];
  assign T2333 = T2338 | T2334;
  assign T2334 = T2335[4'hf:1'h0];
  assign T2335 = T2337 | T2336;
  assign T2336 = hits[5'h1f:1'h0];
  assign T2337 = hits[6'h3d:6'h20];
  assign T2338 = T2335[5'h1f:5'h10];
  assign T2339 = T2333[4'hf:4'h8];
  assign T2340 = T2331[3'h7:3'h4];
  assign T2341 = T2329[2'h3:2'h2];
  assign T2342 = T2341 != 2'h0;
  assign T2343 = T2340 != 4'h0;
  assign T2344 = T2339 != 8'h0;
  assign T2345 = T2338 != 16'h0;
  assign T2346 = T2337 != 30'h0;
  assign io_resp_bits_target = T1406;
  assign T1406 = T2278 ? io_ras_update_bits_returnAddr : T1407;
  assign T1407 = T1900 ? T1867 : T1408;
  assign T1408 = {T1659, T1409};
  assign T1409 = T1416 | T1410;
  assign T1410 = T1415 ? T1411 : 12'h0;
  assign T1411 = tgts[6'h3d];
  assign T2347 = io_req_bits_addr[4'hb:1'h0];
  assign T1413 = R7 & T1414;
  assign T1414 = T42 < 6'h3e;
  assign T1415 = hits[6'h3d:6'h3d];
  assign T1416 = T1420 | T1417;
  assign T1417 = T1419 ? T1418 : 12'h0;
  assign T1418 = tgts[6'h3c];
  assign T1419 = hits[6'h3c:6'h3c];
  assign T1420 = T1424 | T1421;
  assign T1421 = T1423 ? T1422 : 12'h0;
  assign T1422 = tgts[6'h3b];
  assign T1423 = hits[6'h3b:6'h3b];
  assign T1424 = T1428 | T1425;
  assign T1425 = T1427 ? T1426 : 12'h0;
  assign T1426 = tgts[6'h3a];
  assign T1427 = hits[6'h3a:6'h3a];
  assign T1428 = T1432 | T1429;
  assign T1429 = T1431 ? T1430 : 12'h0;
  assign T1430 = tgts[6'h39];
  assign T1431 = hits[6'h39:6'h39];
  assign T1432 = T1436 | T1433;
  assign T1433 = T1435 ? T1434 : 12'h0;
  assign T1434 = tgts[6'h38];
  assign T1435 = hits[6'h38:6'h38];
  assign T1436 = T1440 | T1437;
  assign T1437 = T1439 ? T1438 : 12'h0;
  assign T1438 = tgts[6'h37];
  assign T1439 = hits[6'h37:6'h37];
  assign T1440 = T1444 | T1441;
  assign T1441 = T1443 ? T1442 : 12'h0;
  assign T1442 = tgts[6'h36];
  assign T1443 = hits[6'h36:6'h36];
  assign T1444 = T1448 | T1445;
  assign T1445 = T1447 ? T1446 : 12'h0;
  assign T1446 = tgts[6'h35];
  assign T1447 = hits[6'h35:6'h35];
  assign T1448 = T1452 | T1449;
  assign T1449 = T1451 ? T1450 : 12'h0;
  assign T1450 = tgts[6'h34];
  assign T1451 = hits[6'h34:6'h34];
  assign T1452 = T1456 | T1453;
  assign T1453 = T1455 ? T1454 : 12'h0;
  assign T1454 = tgts[6'h33];
  assign T1455 = hits[6'h33:6'h33];
  assign T1456 = T1460 | T1457;
  assign T1457 = T1459 ? T1458 : 12'h0;
  assign T1458 = tgts[6'h32];
  assign T1459 = hits[6'h32:6'h32];
  assign T1460 = T1464 | T1461;
  assign T1461 = T1463 ? T1462 : 12'h0;
  assign T1462 = tgts[6'h31];
  assign T1463 = hits[6'h31:6'h31];
  assign T1464 = T1468 | T1465;
  assign T1465 = T1467 ? T1466 : 12'h0;
  assign T1466 = tgts[6'h30];
  assign T1467 = hits[6'h30:6'h30];
  assign T1468 = T1472 | T1469;
  assign T1469 = T1471 ? T1470 : 12'h0;
  assign T1470 = tgts[6'h2f];
  assign T1471 = hits[6'h2f:6'h2f];
  assign T1472 = T1476 | T1473;
  assign T1473 = T1475 ? T1474 : 12'h0;
  assign T1474 = tgts[6'h2e];
  assign T1475 = hits[6'h2e:6'h2e];
  assign T1476 = T1480 | T1477;
  assign T1477 = T1479 ? T1478 : 12'h0;
  assign T1478 = tgts[6'h2d];
  assign T1479 = hits[6'h2d:6'h2d];
  assign T1480 = T1484 | T1481;
  assign T1481 = T1483 ? T1482 : 12'h0;
  assign T1482 = tgts[6'h2c];
  assign T1483 = hits[6'h2c:6'h2c];
  assign T1484 = T1488 | T1485;
  assign T1485 = T1487 ? T1486 : 12'h0;
  assign T1486 = tgts[6'h2b];
  assign T1487 = hits[6'h2b:6'h2b];
  assign T1488 = T1492 | T1489;
  assign T1489 = T1491 ? T1490 : 12'h0;
  assign T1490 = tgts[6'h2a];
  assign T1491 = hits[6'h2a:6'h2a];
  assign T1492 = T1496 | T1493;
  assign T1493 = T1495 ? T1494 : 12'h0;
  assign T1494 = tgts[6'h29];
  assign T1495 = hits[6'h29:6'h29];
  assign T1496 = T1500 | T1497;
  assign T1497 = T1499 ? T1498 : 12'h0;
  assign T1498 = tgts[6'h28];
  assign T1499 = hits[6'h28:6'h28];
  assign T1500 = T1504 | T1501;
  assign T1501 = T1503 ? T1502 : 12'h0;
  assign T1502 = tgts[6'h27];
  assign T1503 = hits[6'h27:6'h27];
  assign T1504 = T1508 | T1505;
  assign T1505 = T1507 ? T1506 : 12'h0;
  assign T1506 = tgts[6'h26];
  assign T1507 = hits[6'h26:6'h26];
  assign T1508 = T1512 | T1509;
  assign T1509 = T1511 ? T1510 : 12'h0;
  assign T1510 = tgts[6'h25];
  assign T1511 = hits[6'h25:6'h25];
  assign T1512 = T1516 | T1513;
  assign T1513 = T1515 ? T1514 : 12'h0;
  assign T1514 = tgts[6'h24];
  assign T1515 = hits[6'h24:6'h24];
  assign T1516 = T1520 | T1517;
  assign T1517 = T1519 ? T1518 : 12'h0;
  assign T1518 = tgts[6'h23];
  assign T1519 = hits[6'h23:6'h23];
  assign T1520 = T1524 | T1521;
  assign T1521 = T1523 ? T1522 : 12'h0;
  assign T1522 = tgts[6'h22];
  assign T1523 = hits[6'h22:6'h22];
  assign T1524 = T1528 | T1525;
  assign T1525 = T1527 ? T1526 : 12'h0;
  assign T1526 = tgts[6'h21];
  assign T1527 = hits[6'h21:6'h21];
  assign T1528 = T1532 | T1529;
  assign T1529 = T1531 ? T1530 : 12'h0;
  assign T1530 = tgts[6'h20];
  assign T1531 = hits[6'h20:6'h20];
  assign T1532 = T1536 | T1533;
  assign T1533 = T1535 ? T1534 : 12'h0;
  assign T1534 = tgts[6'h1f];
  assign T1535 = hits[5'h1f:5'h1f];
  assign T1536 = T1540 | T1537;
  assign T1537 = T1539 ? T1538 : 12'h0;
  assign T1538 = tgts[6'h1e];
  assign T1539 = hits[5'h1e:5'h1e];
  assign T1540 = T1544 | T1541;
  assign T1541 = T1543 ? T1542 : 12'h0;
  assign T1542 = tgts[6'h1d];
  assign T1543 = hits[5'h1d:5'h1d];
  assign T1544 = T1548 | T1545;
  assign T1545 = T1547 ? T1546 : 12'h0;
  assign T1546 = tgts[6'h1c];
  assign T1547 = hits[5'h1c:5'h1c];
  assign T1548 = T1552 | T1549;
  assign T1549 = T1551 ? T1550 : 12'h0;
  assign T1550 = tgts[6'h1b];
  assign T1551 = hits[5'h1b:5'h1b];
  assign T1552 = T1556 | T1553;
  assign T1553 = T1555 ? T1554 : 12'h0;
  assign T1554 = tgts[6'h1a];
  assign T1555 = hits[5'h1a:5'h1a];
  assign T1556 = T1560 | T1557;
  assign T1557 = T1559 ? T1558 : 12'h0;
  assign T1558 = tgts[6'h19];
  assign T1559 = hits[5'h19:5'h19];
  assign T1560 = T1564 | T1561;
  assign T1561 = T1563 ? T1562 : 12'h0;
  assign T1562 = tgts[6'h18];
  assign T1563 = hits[5'h18:5'h18];
  assign T1564 = T1568 | T1565;
  assign T1565 = T1567 ? T1566 : 12'h0;
  assign T1566 = tgts[6'h17];
  assign T1567 = hits[5'h17:5'h17];
  assign T1568 = T1572 | T1569;
  assign T1569 = T1571 ? T1570 : 12'h0;
  assign T1570 = tgts[6'h16];
  assign T1571 = hits[5'h16:5'h16];
  assign T1572 = T1576 | T1573;
  assign T1573 = T1575 ? T1574 : 12'h0;
  assign T1574 = tgts[6'h15];
  assign T1575 = hits[5'h15:5'h15];
  assign T1576 = T1580 | T1577;
  assign T1577 = T1579 ? T1578 : 12'h0;
  assign T1578 = tgts[6'h14];
  assign T1579 = hits[5'h14:5'h14];
  assign T1580 = T1584 | T1581;
  assign T1581 = T1583 ? T1582 : 12'h0;
  assign T1582 = tgts[6'h13];
  assign T1583 = hits[5'h13:5'h13];
  assign T1584 = T1588 | T1585;
  assign T1585 = T1587 ? T1586 : 12'h0;
  assign T1586 = tgts[6'h12];
  assign T1587 = hits[5'h12:5'h12];
  assign T1588 = T1592 | T1589;
  assign T1589 = T1591 ? T1590 : 12'h0;
  assign T1590 = tgts[6'h11];
  assign T1591 = hits[5'h11:5'h11];
  assign T1592 = T1596 | T1593;
  assign T1593 = T1595 ? T1594 : 12'h0;
  assign T1594 = tgts[6'h10];
  assign T1595 = hits[5'h10:5'h10];
  assign T1596 = T1600 | T1597;
  assign T1597 = T1599 ? T1598 : 12'h0;
  assign T1598 = tgts[6'hf];
  assign T1599 = hits[4'hf:4'hf];
  assign T1600 = T1604 | T1601;
  assign T1601 = T1603 ? T1602 : 12'h0;
  assign T1602 = tgts[6'he];
  assign T1603 = hits[4'he:4'he];
  assign T1604 = T1608 | T1605;
  assign T1605 = T1607 ? T1606 : 12'h0;
  assign T1606 = tgts[6'hd];
  assign T1607 = hits[4'hd:4'hd];
  assign T1608 = T1612 | T1609;
  assign T1609 = T1611 ? T1610 : 12'h0;
  assign T1610 = tgts[6'hc];
  assign T1611 = hits[4'hc:4'hc];
  assign T1612 = T1616 | T1613;
  assign T1613 = T1615 ? T1614 : 12'h0;
  assign T1614 = tgts[6'hb];
  assign T1615 = hits[4'hb:4'hb];
  assign T1616 = T1620 | T1617;
  assign T1617 = T1619 ? T1618 : 12'h0;
  assign T1618 = tgts[6'ha];
  assign T1619 = hits[4'ha:4'ha];
  assign T1620 = T1624 | T1621;
  assign T1621 = T1623 ? T1622 : 12'h0;
  assign T1622 = tgts[6'h9];
  assign T1623 = hits[4'h9:4'h9];
  assign T1624 = T1628 | T1625;
  assign T1625 = T1627 ? T1626 : 12'h0;
  assign T1626 = tgts[6'h8];
  assign T1627 = hits[4'h8:4'h8];
  assign T1628 = T1632 | T1629;
  assign T1629 = T1631 ? T1630 : 12'h0;
  assign T1630 = tgts[6'h7];
  assign T1631 = hits[3'h7:3'h7];
  assign T1632 = T1636 | T1633;
  assign T1633 = T1635 ? T1634 : 12'h0;
  assign T1634 = tgts[6'h6];
  assign T1635 = hits[3'h6:3'h6];
  assign T1636 = T1640 | T1637;
  assign T1637 = T1639 ? T1638 : 12'h0;
  assign T1638 = tgts[6'h5];
  assign T1639 = hits[3'h5:3'h5];
  assign T1640 = T1644 | T1641;
  assign T1641 = T1643 ? T1642 : 12'h0;
  assign T1642 = tgts[6'h4];
  assign T1643 = hits[3'h4:3'h4];
  assign T1644 = T1648 | T1645;
  assign T1645 = T1647 ? T1646 : 12'h0;
  assign T1646 = tgts[6'h3];
  assign T1647 = hits[2'h3:2'h3];
  assign T1648 = T1652 | T1649;
  assign T1649 = T1651 ? T1650 : 12'h0;
  assign T1650 = tgts[6'h2];
  assign T1651 = hits[2'h2:2'h2];
  assign T1652 = T1656 | T1653;
  assign T1653 = T1655 ? T1654 : 12'h0;
  assign T1654 = tgts[6'h1];
  assign T1655 = hits[1'h1:1'h1];
  assign T1656 = T1658 ? T1657 : 12'h0;
  assign T1657 = tgts[6'h0];
  assign T1658 = hits[1'h0:1'h0];
  assign T1659 = T1848 | T1660;
  assign T1660 = T1662 ? T1661 : 27'h0;
  assign T1661 = pages[3'h5];
  assign T1662 = T1663[3'h5:3'h5];
  assign T1663 = T1666 | T1664;
  assign T1664 = T1665 ? tgtPagesOH_61 : 6'h0;
  assign T1665 = hits[6'h3d:6'h3d];
  assign T1666 = T1669 | T1667;
  assign T1667 = T1668 ? tgtPagesOH_60 : 6'h0;
  assign T1668 = hits[6'h3c:6'h3c];
  assign T1669 = T1672 | T1670;
  assign T1670 = T1671 ? tgtPagesOH_59 : 6'h0;
  assign T1671 = hits[6'h3b:6'h3b];
  assign T1672 = T1675 | T1673;
  assign T1673 = T1674 ? tgtPagesOH_58 : 6'h0;
  assign T1674 = hits[6'h3a:6'h3a];
  assign T1675 = T1678 | T1676;
  assign T1676 = T1677 ? tgtPagesOH_57 : 6'h0;
  assign T1677 = hits[6'h39:6'h39];
  assign T1678 = T1681 | T1679;
  assign T1679 = T1680 ? tgtPagesOH_56 : 6'h0;
  assign T1680 = hits[6'h38:6'h38];
  assign T1681 = T1684 | T1682;
  assign T1682 = T1683 ? tgtPagesOH_55 : 6'h0;
  assign T1683 = hits[6'h37:6'h37];
  assign T1684 = T1687 | T1685;
  assign T1685 = T1686 ? tgtPagesOH_54 : 6'h0;
  assign T1686 = hits[6'h36:6'h36];
  assign T1687 = T1690 | T1688;
  assign T1688 = T1689 ? tgtPagesOH_53 : 6'h0;
  assign T1689 = hits[6'h35:6'h35];
  assign T1690 = T1693 | T1691;
  assign T1691 = T1692 ? tgtPagesOH_52 : 6'h0;
  assign T1692 = hits[6'h34:6'h34];
  assign T1693 = T1696 | T1694;
  assign T1694 = T1695 ? tgtPagesOH_51 : 6'h0;
  assign T1695 = hits[6'h33:6'h33];
  assign T1696 = T1699 | T1697;
  assign T1697 = T1698 ? tgtPagesOH_50 : 6'h0;
  assign T1698 = hits[6'h32:6'h32];
  assign T1699 = T1702 | T1700;
  assign T1700 = T1701 ? tgtPagesOH_49 : 6'h0;
  assign T1701 = hits[6'h31:6'h31];
  assign T1702 = T1705 | T1703;
  assign T1703 = T1704 ? tgtPagesOH_48 : 6'h0;
  assign T1704 = hits[6'h30:6'h30];
  assign T1705 = T1708 | T1706;
  assign T1706 = T1707 ? tgtPagesOH_47 : 6'h0;
  assign T1707 = hits[6'h2f:6'h2f];
  assign T1708 = T1711 | T1709;
  assign T1709 = T1710 ? tgtPagesOH_46 : 6'h0;
  assign T1710 = hits[6'h2e:6'h2e];
  assign T1711 = T1714 | T1712;
  assign T1712 = T1713 ? tgtPagesOH_45 : 6'h0;
  assign T1713 = hits[6'h2d:6'h2d];
  assign T1714 = T1717 | T1715;
  assign T1715 = T1716 ? tgtPagesOH_44 : 6'h0;
  assign T1716 = hits[6'h2c:6'h2c];
  assign T1717 = T1720 | T1718;
  assign T1718 = T1719 ? tgtPagesOH_43 : 6'h0;
  assign T1719 = hits[6'h2b:6'h2b];
  assign T1720 = T1723 | T1721;
  assign T1721 = T1722 ? tgtPagesOH_42 : 6'h0;
  assign T1722 = hits[6'h2a:6'h2a];
  assign T1723 = T1726 | T1724;
  assign T1724 = T1725 ? tgtPagesOH_41 : 6'h0;
  assign T1725 = hits[6'h29:6'h29];
  assign T1726 = T1729 | T1727;
  assign T1727 = T1728 ? tgtPagesOH_40 : 6'h0;
  assign T1728 = hits[6'h28:6'h28];
  assign T1729 = T1732 | T1730;
  assign T1730 = T1731 ? tgtPagesOH_39 : 6'h0;
  assign T1731 = hits[6'h27:6'h27];
  assign T1732 = T1735 | T1733;
  assign T1733 = T1734 ? tgtPagesOH_38 : 6'h0;
  assign T1734 = hits[6'h26:6'h26];
  assign T1735 = T1738 | T1736;
  assign T1736 = T1737 ? tgtPagesOH_37 : 6'h0;
  assign T1737 = hits[6'h25:6'h25];
  assign T1738 = T1741 | T1739;
  assign T1739 = T1740 ? tgtPagesOH_36 : 6'h0;
  assign T1740 = hits[6'h24:6'h24];
  assign T1741 = T1744 | T1742;
  assign T1742 = T1743 ? tgtPagesOH_35 : 6'h0;
  assign T1743 = hits[6'h23:6'h23];
  assign T1744 = T1747 | T1745;
  assign T1745 = T1746 ? tgtPagesOH_34 : 6'h0;
  assign T1746 = hits[6'h22:6'h22];
  assign T1747 = T1750 | T1748;
  assign T1748 = T1749 ? tgtPagesOH_33 : 6'h0;
  assign T1749 = hits[6'h21:6'h21];
  assign T1750 = T1753 | T1751;
  assign T1751 = T1752 ? tgtPagesOH_32 : 6'h0;
  assign T1752 = hits[6'h20:6'h20];
  assign T1753 = T1756 | T1754;
  assign T1754 = T1755 ? tgtPagesOH_31 : 6'h0;
  assign T1755 = hits[5'h1f:5'h1f];
  assign T1756 = T1759 | T1757;
  assign T1757 = T1758 ? tgtPagesOH_30 : 6'h0;
  assign T1758 = hits[5'h1e:5'h1e];
  assign T1759 = T1762 | T1760;
  assign T1760 = T1761 ? tgtPagesOH_29 : 6'h0;
  assign T1761 = hits[5'h1d:5'h1d];
  assign T1762 = T1765 | T1763;
  assign T1763 = T1764 ? tgtPagesOH_28 : 6'h0;
  assign T1764 = hits[5'h1c:5'h1c];
  assign T1765 = T1768 | T1766;
  assign T1766 = T1767 ? tgtPagesOH_27 : 6'h0;
  assign T1767 = hits[5'h1b:5'h1b];
  assign T1768 = T1771 | T1769;
  assign T1769 = T1770 ? tgtPagesOH_26 : 6'h0;
  assign T1770 = hits[5'h1a:5'h1a];
  assign T1771 = T1774 | T1772;
  assign T1772 = T1773 ? tgtPagesOH_25 : 6'h0;
  assign T1773 = hits[5'h19:5'h19];
  assign T1774 = T1777 | T1775;
  assign T1775 = T1776 ? tgtPagesOH_24 : 6'h0;
  assign T1776 = hits[5'h18:5'h18];
  assign T1777 = T1780 | T1778;
  assign T1778 = T1779 ? tgtPagesOH_23 : 6'h0;
  assign T1779 = hits[5'h17:5'h17];
  assign T1780 = T1783 | T1781;
  assign T1781 = T1782 ? tgtPagesOH_22 : 6'h0;
  assign T1782 = hits[5'h16:5'h16];
  assign T1783 = T1786 | T1784;
  assign T1784 = T1785 ? tgtPagesOH_21 : 6'h0;
  assign T1785 = hits[5'h15:5'h15];
  assign T1786 = T1789 | T1787;
  assign T1787 = T1788 ? tgtPagesOH_20 : 6'h0;
  assign T1788 = hits[5'h14:5'h14];
  assign T1789 = T1792 | T1790;
  assign T1790 = T1791 ? tgtPagesOH_19 : 6'h0;
  assign T1791 = hits[5'h13:5'h13];
  assign T1792 = T1795 | T1793;
  assign T1793 = T1794 ? tgtPagesOH_18 : 6'h0;
  assign T1794 = hits[5'h12:5'h12];
  assign T1795 = T1798 | T1796;
  assign T1796 = T1797 ? tgtPagesOH_17 : 6'h0;
  assign T1797 = hits[5'h11:5'h11];
  assign T1798 = T1801 | T1799;
  assign T1799 = T1800 ? tgtPagesOH_16 : 6'h0;
  assign T1800 = hits[5'h10:5'h10];
  assign T1801 = T1804 | T1802;
  assign T1802 = T1803 ? tgtPagesOH_15 : 6'h0;
  assign T1803 = hits[4'hf:4'hf];
  assign T1804 = T1807 | T1805;
  assign T1805 = T1806 ? tgtPagesOH_14 : 6'h0;
  assign T1806 = hits[4'he:4'he];
  assign T1807 = T1810 | T1808;
  assign T1808 = T1809 ? tgtPagesOH_13 : 6'h0;
  assign T1809 = hits[4'hd:4'hd];
  assign T1810 = T1813 | T1811;
  assign T1811 = T1812 ? tgtPagesOH_12 : 6'h0;
  assign T1812 = hits[4'hc:4'hc];
  assign T1813 = T1816 | T1814;
  assign T1814 = T1815 ? tgtPagesOH_11 : 6'h0;
  assign T1815 = hits[4'hb:4'hb];
  assign T1816 = T1819 | T1817;
  assign T1817 = T1818 ? tgtPagesOH_10 : 6'h0;
  assign T1818 = hits[4'ha:4'ha];
  assign T1819 = T1822 | T1820;
  assign T1820 = T1821 ? tgtPagesOH_9 : 6'h0;
  assign T1821 = hits[4'h9:4'h9];
  assign T1822 = T1825 | T1823;
  assign T1823 = T1824 ? tgtPagesOH_8 : 6'h0;
  assign T1824 = hits[4'h8:4'h8];
  assign T1825 = T1828 | T1826;
  assign T1826 = T1827 ? tgtPagesOH_7 : 6'h0;
  assign T1827 = hits[3'h7:3'h7];
  assign T1828 = T1831 | T1829;
  assign T1829 = T1830 ? tgtPagesOH_6 : 6'h0;
  assign T1830 = hits[3'h6:3'h6];
  assign T1831 = T1834 | T1832;
  assign T1832 = T1833 ? tgtPagesOH_5 : 6'h0;
  assign T1833 = hits[3'h5:3'h5];
  assign T1834 = T1837 | T1835;
  assign T1835 = T1836 ? tgtPagesOH_4 : 6'h0;
  assign T1836 = hits[3'h4:3'h4];
  assign T1837 = T1840 | T1838;
  assign T1838 = T1839 ? tgtPagesOH_3 : 6'h0;
  assign T1839 = hits[2'h3:2'h3];
  assign T1840 = T1843 | T1841;
  assign T1841 = T1842 ? tgtPagesOH_2 : 6'h0;
  assign T1842 = hits[2'h2:2'h2];
  assign T1843 = T1846 | T1844;
  assign T1844 = T1845 ? tgtPagesOH_1 : 6'h0;
  assign T1845 = hits[1'h1:1'h1];
  assign T1846 = T1847 ? tgtPagesOH_0 : 6'h0;
  assign T1847 = hits[1'h0:1'h0];
  assign T1848 = T1852 | T1849;
  assign T1849 = T1851 ? T1850 : 27'h0;
  assign T1850 = pages[3'h4];
  assign T1851 = T1663[3'h4:3'h4];
  assign T1852 = T1856 | T1853;
  assign T1853 = T1855 ? T1854 : 27'h0;
  assign T1854 = pages[3'h3];
  assign T1855 = T1663[2'h3:2'h3];
  assign T1856 = T1860 | T1857;
  assign T1857 = T1859 ? T1858 : 27'h0;
  assign T1858 = pages[3'h2];
  assign T1859 = T1663[2'h2:2'h2];
  assign T1860 = T1864 | T1861;
  assign T1861 = T1863 ? T1862 : 27'h0;
  assign T1862 = pages[3'h1];
  assign T1863 = T1663[1'h1:1'h1];
  assign T1864 = T1866 ? T1865 : 27'h0;
  assign T1865 = pages[3'h0];
  assign T1866 = T1663[1'h0:1'h0];
  assign T1867 = T1899 ? R1895 : R1868;
  assign T1869 = T1870 ? io_ras_update_bits_returnAddr : R1868;
  assign T1870 = T1894 & T1871;
  assign T1871 = T1872[1'h0:1'h0];
  assign T1872 = 1'h1 << T1873;
  assign T1873 = T1874;
  assign T1874 = R1875 + 1'h1;
  assign T2348 = reset ? 1'h0 : T1876;
  assign T1876 = T1879 ? T1878 : T1877;
  assign T1877 = T1894 ? T1874 : R1875;
  assign T1878 = R1875 - 1'h1;
  assign T1879 = T1890 & T1880;
  assign T1880 = T1881 ^ 1'h1;
  assign T1881 = R1882 == 2'h0;
  assign T2349 = reset ? 2'h0 : T1883;
  assign T1883 = io_invalidate ? 2'h0 : T1884;
  assign T1884 = T1879 ? T1889 : T1885;
  assign T1885 = T1887 ? T1886 : R1882;
  assign T1886 = R1882 + 2'h1;
  assign T1887 = T1894 & T1888;
  assign T1888 = R1882 < 2'h2;
  assign T1889 = R1882 - 2'h1;
  assign T1890 = io_ras_update_valid & T1891;
  assign T1891 = T1893 & T1892;
  assign T1892 = io_ras_update_bits_isReturn & io_ras_update_bits_prediction_valid;
  assign T1893 = io_ras_update_bits_isCall ^ 1'h1;
  assign T1894 = io_ras_update_valid & io_ras_update_bits_isCall;
  assign T1896 = T1897 ? io_ras_update_bits_returnAddr : R1895;
  assign T1897 = T1894 & T1898;
  assign T1898 = T1872[1'h1:1'h1];
  assign T1899 = R1875;
  assign T1900 = T2276 & T1901;
  assign T1901 = T1911 | T1902;
  assign T1902 = T1910 ? useRAS_61 : 1'h0;
  assign T1903 = T1906 ? R1904 : useRAS_61;
  assign T1905 = io_btb_update_valid ? io_btb_update_bits_isReturn : R1904;
  assign T1906 = R7 & T1907;
  assign T1907 = T1908[6'h3d:6'h3d];
  assign T1908 = 1'h1 << T1909;
  assign T1909 = T42;
  assign T1910 = hits[6'h3d:6'h3d];
  assign T1911 = T1917 | T1912;
  assign T1912 = T1916 ? useRAS_60 : 1'h0;
  assign T1913 = T1914 ? R1904 : useRAS_60;
  assign T1914 = R7 & T1915;
  assign T1915 = T1908[6'h3c:6'h3c];
  assign T1916 = hits[6'h3c:6'h3c];
  assign T1917 = T1923 | T1918;
  assign T1918 = T1922 ? useRAS_59 : 1'h0;
  assign T1919 = T1920 ? R1904 : useRAS_59;
  assign T1920 = R7 & T1921;
  assign T1921 = T1908[6'h3b:6'h3b];
  assign T1922 = hits[6'h3b:6'h3b];
  assign T1923 = T1929 | T1924;
  assign T1924 = T1928 ? useRAS_58 : 1'h0;
  assign T1925 = T1926 ? R1904 : useRAS_58;
  assign T1926 = R7 & T1927;
  assign T1927 = T1908[6'h3a:6'h3a];
  assign T1928 = hits[6'h3a:6'h3a];
  assign T1929 = T1935 | T1930;
  assign T1930 = T1934 ? useRAS_57 : 1'h0;
  assign T1931 = T1932 ? R1904 : useRAS_57;
  assign T1932 = R7 & T1933;
  assign T1933 = T1908[6'h39:6'h39];
  assign T1934 = hits[6'h39:6'h39];
  assign T1935 = T1941 | T1936;
  assign T1936 = T1940 ? useRAS_56 : 1'h0;
  assign T1937 = T1938 ? R1904 : useRAS_56;
  assign T1938 = R7 & T1939;
  assign T1939 = T1908[6'h38:6'h38];
  assign T1940 = hits[6'h38:6'h38];
  assign T1941 = T1947 | T1942;
  assign T1942 = T1946 ? useRAS_55 : 1'h0;
  assign T1943 = T1944 ? R1904 : useRAS_55;
  assign T1944 = R7 & T1945;
  assign T1945 = T1908[6'h37:6'h37];
  assign T1946 = hits[6'h37:6'h37];
  assign T1947 = T1953 | T1948;
  assign T1948 = T1952 ? useRAS_54 : 1'h0;
  assign T1949 = T1950 ? R1904 : useRAS_54;
  assign T1950 = R7 & T1951;
  assign T1951 = T1908[6'h36:6'h36];
  assign T1952 = hits[6'h36:6'h36];
  assign T1953 = T1959 | T1954;
  assign T1954 = T1958 ? useRAS_53 : 1'h0;
  assign T1955 = T1956 ? R1904 : useRAS_53;
  assign T1956 = R7 & T1957;
  assign T1957 = T1908[6'h35:6'h35];
  assign T1958 = hits[6'h35:6'h35];
  assign T1959 = T1965 | T1960;
  assign T1960 = T1964 ? useRAS_52 : 1'h0;
  assign T1961 = T1962 ? R1904 : useRAS_52;
  assign T1962 = R7 & T1963;
  assign T1963 = T1908[6'h34:6'h34];
  assign T1964 = hits[6'h34:6'h34];
  assign T1965 = T1971 | T1966;
  assign T1966 = T1970 ? useRAS_51 : 1'h0;
  assign T1967 = T1968 ? R1904 : useRAS_51;
  assign T1968 = R7 & T1969;
  assign T1969 = T1908[6'h33:6'h33];
  assign T1970 = hits[6'h33:6'h33];
  assign T1971 = T1977 | T1972;
  assign T1972 = T1976 ? useRAS_50 : 1'h0;
  assign T1973 = T1974 ? R1904 : useRAS_50;
  assign T1974 = R7 & T1975;
  assign T1975 = T1908[6'h32:6'h32];
  assign T1976 = hits[6'h32:6'h32];
  assign T1977 = T1983 | T1978;
  assign T1978 = T1982 ? useRAS_49 : 1'h0;
  assign T1979 = T1980 ? R1904 : useRAS_49;
  assign T1980 = R7 & T1981;
  assign T1981 = T1908[6'h31:6'h31];
  assign T1982 = hits[6'h31:6'h31];
  assign T1983 = T1989 | T1984;
  assign T1984 = T1988 ? useRAS_48 : 1'h0;
  assign T1985 = T1986 ? R1904 : useRAS_48;
  assign T1986 = R7 & T1987;
  assign T1987 = T1908[6'h30:6'h30];
  assign T1988 = hits[6'h30:6'h30];
  assign T1989 = T1995 | T1990;
  assign T1990 = T1994 ? useRAS_47 : 1'h0;
  assign T1991 = T1992 ? R1904 : useRAS_47;
  assign T1992 = R7 & T1993;
  assign T1993 = T1908[6'h2f:6'h2f];
  assign T1994 = hits[6'h2f:6'h2f];
  assign T1995 = T2001 | T1996;
  assign T1996 = T2000 ? useRAS_46 : 1'h0;
  assign T1997 = T1998 ? R1904 : useRAS_46;
  assign T1998 = R7 & T1999;
  assign T1999 = T1908[6'h2e:6'h2e];
  assign T2000 = hits[6'h2e:6'h2e];
  assign T2001 = T2007 | T2002;
  assign T2002 = T2006 ? useRAS_45 : 1'h0;
  assign T2003 = T2004 ? R1904 : useRAS_45;
  assign T2004 = R7 & T2005;
  assign T2005 = T1908[6'h2d:6'h2d];
  assign T2006 = hits[6'h2d:6'h2d];
  assign T2007 = T2013 | T2008;
  assign T2008 = T2012 ? useRAS_44 : 1'h0;
  assign T2009 = T2010 ? R1904 : useRAS_44;
  assign T2010 = R7 & T2011;
  assign T2011 = T1908[6'h2c:6'h2c];
  assign T2012 = hits[6'h2c:6'h2c];
  assign T2013 = T2019 | T2014;
  assign T2014 = T2018 ? useRAS_43 : 1'h0;
  assign T2015 = T2016 ? R1904 : useRAS_43;
  assign T2016 = R7 & T2017;
  assign T2017 = T1908[6'h2b:6'h2b];
  assign T2018 = hits[6'h2b:6'h2b];
  assign T2019 = T2025 | T2020;
  assign T2020 = T2024 ? useRAS_42 : 1'h0;
  assign T2021 = T2022 ? R1904 : useRAS_42;
  assign T2022 = R7 & T2023;
  assign T2023 = T1908[6'h2a:6'h2a];
  assign T2024 = hits[6'h2a:6'h2a];
  assign T2025 = T2031 | T2026;
  assign T2026 = T2030 ? useRAS_41 : 1'h0;
  assign T2027 = T2028 ? R1904 : useRAS_41;
  assign T2028 = R7 & T2029;
  assign T2029 = T1908[6'h29:6'h29];
  assign T2030 = hits[6'h29:6'h29];
  assign T2031 = T2037 | T2032;
  assign T2032 = T2036 ? useRAS_40 : 1'h0;
  assign T2033 = T2034 ? R1904 : useRAS_40;
  assign T2034 = R7 & T2035;
  assign T2035 = T1908[6'h28:6'h28];
  assign T2036 = hits[6'h28:6'h28];
  assign T2037 = T2043 | T2038;
  assign T2038 = T2042 ? useRAS_39 : 1'h0;
  assign T2039 = T2040 ? R1904 : useRAS_39;
  assign T2040 = R7 & T2041;
  assign T2041 = T1908[6'h27:6'h27];
  assign T2042 = hits[6'h27:6'h27];
  assign T2043 = T2049 | T2044;
  assign T2044 = T2048 ? useRAS_38 : 1'h0;
  assign T2045 = T2046 ? R1904 : useRAS_38;
  assign T2046 = R7 & T2047;
  assign T2047 = T1908[6'h26:6'h26];
  assign T2048 = hits[6'h26:6'h26];
  assign T2049 = T2055 | T2050;
  assign T2050 = T2054 ? useRAS_37 : 1'h0;
  assign T2051 = T2052 ? R1904 : useRAS_37;
  assign T2052 = R7 & T2053;
  assign T2053 = T1908[6'h25:6'h25];
  assign T2054 = hits[6'h25:6'h25];
  assign T2055 = T2061 | T2056;
  assign T2056 = T2060 ? useRAS_36 : 1'h0;
  assign T2057 = T2058 ? R1904 : useRAS_36;
  assign T2058 = R7 & T2059;
  assign T2059 = T1908[6'h24:6'h24];
  assign T2060 = hits[6'h24:6'h24];
  assign T2061 = T2067 | T2062;
  assign T2062 = T2066 ? useRAS_35 : 1'h0;
  assign T2063 = T2064 ? R1904 : useRAS_35;
  assign T2064 = R7 & T2065;
  assign T2065 = T1908[6'h23:6'h23];
  assign T2066 = hits[6'h23:6'h23];
  assign T2067 = T2073 | T2068;
  assign T2068 = T2072 ? useRAS_34 : 1'h0;
  assign T2069 = T2070 ? R1904 : useRAS_34;
  assign T2070 = R7 & T2071;
  assign T2071 = T1908[6'h22:6'h22];
  assign T2072 = hits[6'h22:6'h22];
  assign T2073 = T2079 | T2074;
  assign T2074 = T2078 ? useRAS_33 : 1'h0;
  assign T2075 = T2076 ? R1904 : useRAS_33;
  assign T2076 = R7 & T2077;
  assign T2077 = T1908[6'h21:6'h21];
  assign T2078 = hits[6'h21:6'h21];
  assign T2079 = T2085 | T2080;
  assign T2080 = T2084 ? useRAS_32 : 1'h0;
  assign T2081 = T2082 ? R1904 : useRAS_32;
  assign T2082 = R7 & T2083;
  assign T2083 = T1908[6'h20:6'h20];
  assign T2084 = hits[6'h20:6'h20];
  assign T2085 = T2091 | T2086;
  assign T2086 = T2090 ? useRAS_31 : 1'h0;
  assign T2087 = T2088 ? R1904 : useRAS_31;
  assign T2088 = R7 & T2089;
  assign T2089 = T1908[5'h1f:5'h1f];
  assign T2090 = hits[5'h1f:5'h1f];
  assign T2091 = T2097 | T2092;
  assign T2092 = T2096 ? useRAS_30 : 1'h0;
  assign T2093 = T2094 ? R1904 : useRAS_30;
  assign T2094 = R7 & T2095;
  assign T2095 = T1908[5'h1e:5'h1e];
  assign T2096 = hits[5'h1e:5'h1e];
  assign T2097 = T2103 | T2098;
  assign T2098 = T2102 ? useRAS_29 : 1'h0;
  assign T2099 = T2100 ? R1904 : useRAS_29;
  assign T2100 = R7 & T2101;
  assign T2101 = T1908[5'h1d:5'h1d];
  assign T2102 = hits[5'h1d:5'h1d];
  assign T2103 = T2109 | T2104;
  assign T2104 = T2108 ? useRAS_28 : 1'h0;
  assign T2105 = T2106 ? R1904 : useRAS_28;
  assign T2106 = R7 & T2107;
  assign T2107 = T1908[5'h1c:5'h1c];
  assign T2108 = hits[5'h1c:5'h1c];
  assign T2109 = T2115 | T2110;
  assign T2110 = T2114 ? useRAS_27 : 1'h0;
  assign T2111 = T2112 ? R1904 : useRAS_27;
  assign T2112 = R7 & T2113;
  assign T2113 = T1908[5'h1b:5'h1b];
  assign T2114 = hits[5'h1b:5'h1b];
  assign T2115 = T2121 | T2116;
  assign T2116 = T2120 ? useRAS_26 : 1'h0;
  assign T2117 = T2118 ? R1904 : useRAS_26;
  assign T2118 = R7 & T2119;
  assign T2119 = T1908[5'h1a:5'h1a];
  assign T2120 = hits[5'h1a:5'h1a];
  assign T2121 = T2127 | T2122;
  assign T2122 = T2126 ? useRAS_25 : 1'h0;
  assign T2123 = T2124 ? R1904 : useRAS_25;
  assign T2124 = R7 & T2125;
  assign T2125 = T1908[5'h19:5'h19];
  assign T2126 = hits[5'h19:5'h19];
  assign T2127 = T2133 | T2128;
  assign T2128 = T2132 ? useRAS_24 : 1'h0;
  assign T2129 = T2130 ? R1904 : useRAS_24;
  assign T2130 = R7 & T2131;
  assign T2131 = T1908[5'h18:5'h18];
  assign T2132 = hits[5'h18:5'h18];
  assign T2133 = T2139 | T2134;
  assign T2134 = T2138 ? useRAS_23 : 1'h0;
  assign T2135 = T2136 ? R1904 : useRAS_23;
  assign T2136 = R7 & T2137;
  assign T2137 = T1908[5'h17:5'h17];
  assign T2138 = hits[5'h17:5'h17];
  assign T2139 = T2145 | T2140;
  assign T2140 = T2144 ? useRAS_22 : 1'h0;
  assign T2141 = T2142 ? R1904 : useRAS_22;
  assign T2142 = R7 & T2143;
  assign T2143 = T1908[5'h16:5'h16];
  assign T2144 = hits[5'h16:5'h16];
  assign T2145 = T2151 | T2146;
  assign T2146 = T2150 ? useRAS_21 : 1'h0;
  assign T2147 = T2148 ? R1904 : useRAS_21;
  assign T2148 = R7 & T2149;
  assign T2149 = T1908[5'h15:5'h15];
  assign T2150 = hits[5'h15:5'h15];
  assign T2151 = T2157 | T2152;
  assign T2152 = T2156 ? useRAS_20 : 1'h0;
  assign T2153 = T2154 ? R1904 : useRAS_20;
  assign T2154 = R7 & T2155;
  assign T2155 = T1908[5'h14:5'h14];
  assign T2156 = hits[5'h14:5'h14];
  assign T2157 = T2163 | T2158;
  assign T2158 = T2162 ? useRAS_19 : 1'h0;
  assign T2159 = T2160 ? R1904 : useRAS_19;
  assign T2160 = R7 & T2161;
  assign T2161 = T1908[5'h13:5'h13];
  assign T2162 = hits[5'h13:5'h13];
  assign T2163 = T2169 | T2164;
  assign T2164 = T2168 ? useRAS_18 : 1'h0;
  assign T2165 = T2166 ? R1904 : useRAS_18;
  assign T2166 = R7 & T2167;
  assign T2167 = T1908[5'h12:5'h12];
  assign T2168 = hits[5'h12:5'h12];
  assign T2169 = T2175 | T2170;
  assign T2170 = T2174 ? useRAS_17 : 1'h0;
  assign T2171 = T2172 ? R1904 : useRAS_17;
  assign T2172 = R7 & T2173;
  assign T2173 = T1908[5'h11:5'h11];
  assign T2174 = hits[5'h11:5'h11];
  assign T2175 = T2181 | T2176;
  assign T2176 = T2180 ? useRAS_16 : 1'h0;
  assign T2177 = T2178 ? R1904 : useRAS_16;
  assign T2178 = R7 & T2179;
  assign T2179 = T1908[5'h10:5'h10];
  assign T2180 = hits[5'h10:5'h10];
  assign T2181 = T2187 | T2182;
  assign T2182 = T2186 ? useRAS_15 : 1'h0;
  assign T2183 = T2184 ? R1904 : useRAS_15;
  assign T2184 = R7 & T2185;
  assign T2185 = T1908[4'hf:4'hf];
  assign T2186 = hits[4'hf:4'hf];
  assign T2187 = T2193 | T2188;
  assign T2188 = T2192 ? useRAS_14 : 1'h0;
  assign T2189 = T2190 ? R1904 : useRAS_14;
  assign T2190 = R7 & T2191;
  assign T2191 = T1908[4'he:4'he];
  assign T2192 = hits[4'he:4'he];
  assign T2193 = T2199 | T2194;
  assign T2194 = T2198 ? useRAS_13 : 1'h0;
  assign T2195 = T2196 ? R1904 : useRAS_13;
  assign T2196 = R7 & T2197;
  assign T2197 = T1908[4'hd:4'hd];
  assign T2198 = hits[4'hd:4'hd];
  assign T2199 = T2205 | T2200;
  assign T2200 = T2204 ? useRAS_12 : 1'h0;
  assign T2201 = T2202 ? R1904 : useRAS_12;
  assign T2202 = R7 & T2203;
  assign T2203 = T1908[4'hc:4'hc];
  assign T2204 = hits[4'hc:4'hc];
  assign T2205 = T2211 | T2206;
  assign T2206 = T2210 ? useRAS_11 : 1'h0;
  assign T2207 = T2208 ? R1904 : useRAS_11;
  assign T2208 = R7 & T2209;
  assign T2209 = T1908[4'hb:4'hb];
  assign T2210 = hits[4'hb:4'hb];
  assign T2211 = T2217 | T2212;
  assign T2212 = T2216 ? useRAS_10 : 1'h0;
  assign T2213 = T2214 ? R1904 : useRAS_10;
  assign T2214 = R7 & T2215;
  assign T2215 = T1908[4'ha:4'ha];
  assign T2216 = hits[4'ha:4'ha];
  assign T2217 = T2223 | T2218;
  assign T2218 = T2222 ? useRAS_9 : 1'h0;
  assign T2219 = T2220 ? R1904 : useRAS_9;
  assign T2220 = R7 & T2221;
  assign T2221 = T1908[4'h9:4'h9];
  assign T2222 = hits[4'h9:4'h9];
  assign T2223 = T2229 | T2224;
  assign T2224 = T2228 ? useRAS_8 : 1'h0;
  assign T2225 = T2226 ? R1904 : useRAS_8;
  assign T2226 = R7 & T2227;
  assign T2227 = T1908[4'h8:4'h8];
  assign T2228 = hits[4'h8:4'h8];
  assign T2229 = T2235 | T2230;
  assign T2230 = T2234 ? useRAS_7 : 1'h0;
  assign T2231 = T2232 ? R1904 : useRAS_7;
  assign T2232 = R7 & T2233;
  assign T2233 = T1908[3'h7:3'h7];
  assign T2234 = hits[3'h7:3'h7];
  assign T2235 = T2241 | T2236;
  assign T2236 = T2240 ? useRAS_6 : 1'h0;
  assign T2237 = T2238 ? R1904 : useRAS_6;
  assign T2238 = R7 & T2239;
  assign T2239 = T1908[3'h6:3'h6];
  assign T2240 = hits[3'h6:3'h6];
  assign T2241 = T2247 | T2242;
  assign T2242 = T2246 ? useRAS_5 : 1'h0;
  assign T2243 = T2244 ? R1904 : useRAS_5;
  assign T2244 = R7 & T2245;
  assign T2245 = T1908[3'h5:3'h5];
  assign T2246 = hits[3'h5:3'h5];
  assign T2247 = T2253 | T2248;
  assign T2248 = T2252 ? useRAS_4 : 1'h0;
  assign T2249 = T2250 ? R1904 : useRAS_4;
  assign T2250 = R7 & T2251;
  assign T2251 = T1908[3'h4:3'h4];
  assign T2252 = hits[3'h4:3'h4];
  assign T2253 = T2259 | T2254;
  assign T2254 = T2258 ? useRAS_3 : 1'h0;
  assign T2255 = T2256 ? R1904 : useRAS_3;
  assign T2256 = R7 & T2257;
  assign T2257 = T1908[2'h3:2'h3];
  assign T2258 = hits[2'h3:2'h3];
  assign T2259 = T2265 | T2260;
  assign T2260 = T2264 ? useRAS_2 : 1'h0;
  assign T2261 = T2262 ? R1904 : useRAS_2;
  assign T2262 = R7 & T2263;
  assign T2263 = T1908[2'h2:2'h2];
  assign T2264 = hits[2'h2:2'h2];
  assign T2265 = T2271 | T2266;
  assign T2266 = T2270 ? useRAS_1 : 1'h0;
  assign T2267 = T2268 ? R1904 : useRAS_1;
  assign T2268 = R7 & T2269;
  assign T2269 = T1908[1'h1:1'h1];
  assign T2270 = hits[1'h1:1'h1];
  assign T2271 = T2275 ? useRAS_0 : 1'h0;
  assign T2272 = T2273 ? R1904 : useRAS_0;
  assign T2273 = R7 & T2274;
  assign T2274 = T1908[1'h0:1'h0];
  assign T2275 = hits[1'h0:1'h0];
  assign T2276 = T2277 ^ 1'h1;
  assign T2277 = R1882 == 2'h0;
  assign T2278 = T1894 & T1901;
  assign io_resp_bits_bridx = T2279;
  assign T2279 = brIdx[io_resp_bits_entry];
  assign T2281 = R7 & T2282;
  assign T2282 = T42 < 6'h3e;
  assign io_resp_bits_mask = 1'h1;
  assign io_resp_bits_taken = T2283;
  assign T2283 = T2284 ? 1'h0 : io_resp_valid;
  assign T2284 = T2285 & T32;
  assign T2285 = T2286 ^ 1'h1;
  assign T2286 = T8[1'h0:1'h0];
  assign io_resp_valid = T2287;
  assign T2287 = hits != 62'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
// synthesis translate_on
`endif
    if(io_btb_update_valid) begin
      R4 <= io_btb_update_bits_target;
    end
    if(reset) begin
      R7 <= 1'h0;
    end else begin
      R7 <= io_btb_update_valid;
    end
    if (T21)
      T10[T22] <= T12;
    if(T1402) begin
      R25 <= T1400;
    end else if(T31) begin
      R25 <= T28;
    end
    if(T38) begin
      isJump_61 <= R36;
    end
    if(io_btb_update_valid) begin
      R36 <= io_btb_update_bits_isJump;
    end
    if(reset) begin
      nextRepl <= 6'h0;
    end else if(T47) begin
      nextRepl <= T44;
    end
    if(io_btb_update_valid) begin
      R49 <= io_btb_update_bits_prediction_bits_entry;
    end
    if(io_btb_update_valid) begin
      updateHit <= io_btb_update_bits_prediction_valid;
    end
    if(reset) begin
      pageValid <= 6'h0;
    end else if(io_invalidate) begin
      pageValid <= 6'h0;
    end else if(T137) begin
      pageValid <= T64;
    end
    if(reset) begin
      R70 <= 3'h0;
    end else if(T75) begin
      R70 <= T72;
    end
    if(io_btb_update_valid) begin
      R82 <= io_btb_update_bits_pc;
    end
    if (T91)
      pages[3'h5] <= T86;
    if (T96)
      pages[3'h3] <= T86;
    if (T100)
      pages[3'h1] <= T86;
    if (T107)
      pages[3'h4] <= T104;
    if (T112)
      pages[3'h2] <= T104;
    if (T116)
      pages[3'h0] <= T104;
    if (T160)
      idxPages[T42] <= T2294;
    if (T473)
      idxs[T42] <= T2305;
    idxValid <= T2306;
    if (T672)
      tgtPages[T42] <= T2310;
    if(T1037) begin
      isJump_60 <= R36;
    end
    if(T1043) begin
      isJump_59 <= R36;
    end
    if(T1049) begin
      isJump_58 <= R36;
    end
    if(T1055) begin
      isJump_57 <= R36;
    end
    if(T1061) begin
      isJump_56 <= R36;
    end
    if(T1067) begin
      isJump_55 <= R36;
    end
    if(T1073) begin
      isJump_54 <= R36;
    end
    if(T1079) begin
      isJump_53 <= R36;
    end
    if(T1085) begin
      isJump_52 <= R36;
    end
    if(T1091) begin
      isJump_51 <= R36;
    end
    if(T1097) begin
      isJump_50 <= R36;
    end
    if(T1103) begin
      isJump_49 <= R36;
    end
    if(T1109) begin
      isJump_48 <= R36;
    end
    if(T1115) begin
      isJump_47 <= R36;
    end
    if(T1121) begin
      isJump_46 <= R36;
    end
    if(T1127) begin
      isJump_45 <= R36;
    end
    if(T1133) begin
      isJump_44 <= R36;
    end
    if(T1139) begin
      isJump_43 <= R36;
    end
    if(T1145) begin
      isJump_42 <= R36;
    end
    if(T1151) begin
      isJump_41 <= R36;
    end
    if(T1157) begin
      isJump_40 <= R36;
    end
    if(T1163) begin
      isJump_39 <= R36;
    end
    if(T1169) begin
      isJump_38 <= R36;
    end
    if(T1175) begin
      isJump_37 <= R36;
    end
    if(T1181) begin
      isJump_36 <= R36;
    end
    if(T1187) begin
      isJump_35 <= R36;
    end
    if(T1193) begin
      isJump_34 <= R36;
    end
    if(T1199) begin
      isJump_33 <= R36;
    end
    if(T1205) begin
      isJump_32 <= R36;
    end
    if(T1211) begin
      isJump_31 <= R36;
    end
    if(T1217) begin
      isJump_30 <= R36;
    end
    if(T1223) begin
      isJump_29 <= R36;
    end
    if(T1229) begin
      isJump_28 <= R36;
    end
    if(T1235) begin
      isJump_27 <= R36;
    end
    if(T1241) begin
      isJump_26 <= R36;
    end
    if(T1247) begin
      isJump_25 <= R36;
    end
    if(T1253) begin
      isJump_24 <= R36;
    end
    if(T1259) begin
      isJump_23 <= R36;
    end
    if(T1265) begin
      isJump_22 <= R36;
    end
    if(T1271) begin
      isJump_21 <= R36;
    end
    if(T1277) begin
      isJump_20 <= R36;
    end
    if(T1283) begin
      isJump_19 <= R36;
    end
    if(T1289) begin
      isJump_18 <= R36;
    end
    if(T1295) begin
      isJump_17 <= R36;
    end
    if(T1301) begin
      isJump_16 <= R36;
    end
    if(T1307) begin
      isJump_15 <= R36;
    end
    if(T1313) begin
      isJump_14 <= R36;
    end
    if(T1319) begin
      isJump_13 <= R36;
    end
    if(T1325) begin
      isJump_12 <= R36;
    end
    if(T1331) begin
      isJump_11 <= R36;
    end
    if(T1337) begin
      isJump_10 <= R36;
    end
    if(T1343) begin
      isJump_9 <= R36;
    end
    if(T1349) begin
      isJump_8 <= R36;
    end
    if(T1355) begin
      isJump_7 <= R36;
    end
    if(T1361) begin
      isJump_6 <= R36;
    end
    if(T1367) begin
      isJump_5 <= R36;
    end
    if(T1373) begin
      isJump_4 <= R36;
    end
    if(T1379) begin
      isJump_3 <= R36;
    end
    if(T1385) begin
      isJump_2 <= R36;
    end
    if(T1391) begin
      isJump_1 <= R36;
    end
    if(T1396) begin
      isJump_0 <= R36;
    end
    if (T1413)
      tgts[T42] <= T2347;
    if(T1870) begin
      R1868 <= io_ras_update_bits_returnAddr;
    end
    if(reset) begin
      R1875 <= 1'h0;
    end else if(T1879) begin
      R1875 <= T1878;
    end else if(T1894) begin
      R1875 <= T1874;
    end
    if(reset) begin
      R1882 <= 2'h0;
    end else if(io_invalidate) begin
      R1882 <= 2'h0;
    end else if(T1879) begin
      R1882 <= T1889;
    end else if(T1887) begin
      R1882 <= T1886;
    end
    if(T1897) begin
      R1895 <= io_ras_update_bits_returnAddr;
    end
    if(T1906) begin
      useRAS_61 <= R1904;
    end
    if(io_btb_update_valid) begin
      R1904 <= io_btb_update_bits_isReturn;
    end
    if(T1914) begin
      useRAS_60 <= R1904;
    end
    if(T1920) begin
      useRAS_59 <= R1904;
    end
    if(T1926) begin
      useRAS_58 <= R1904;
    end
    if(T1932) begin
      useRAS_57 <= R1904;
    end
    if(T1938) begin
      useRAS_56 <= R1904;
    end
    if(T1944) begin
      useRAS_55 <= R1904;
    end
    if(T1950) begin
      useRAS_54 <= R1904;
    end
    if(T1956) begin
      useRAS_53 <= R1904;
    end
    if(T1962) begin
      useRAS_52 <= R1904;
    end
    if(T1968) begin
      useRAS_51 <= R1904;
    end
    if(T1974) begin
      useRAS_50 <= R1904;
    end
    if(T1980) begin
      useRAS_49 <= R1904;
    end
    if(T1986) begin
      useRAS_48 <= R1904;
    end
    if(T1992) begin
      useRAS_47 <= R1904;
    end
    if(T1998) begin
      useRAS_46 <= R1904;
    end
    if(T2004) begin
      useRAS_45 <= R1904;
    end
    if(T2010) begin
      useRAS_44 <= R1904;
    end
    if(T2016) begin
      useRAS_43 <= R1904;
    end
    if(T2022) begin
      useRAS_42 <= R1904;
    end
    if(T2028) begin
      useRAS_41 <= R1904;
    end
    if(T2034) begin
      useRAS_40 <= R1904;
    end
    if(T2040) begin
      useRAS_39 <= R1904;
    end
    if(T2046) begin
      useRAS_38 <= R1904;
    end
    if(T2052) begin
      useRAS_37 <= R1904;
    end
    if(T2058) begin
      useRAS_36 <= R1904;
    end
    if(T2064) begin
      useRAS_35 <= R1904;
    end
    if(T2070) begin
      useRAS_34 <= R1904;
    end
    if(T2076) begin
      useRAS_33 <= R1904;
    end
    if(T2082) begin
      useRAS_32 <= R1904;
    end
    if(T2088) begin
      useRAS_31 <= R1904;
    end
    if(T2094) begin
      useRAS_30 <= R1904;
    end
    if(T2100) begin
      useRAS_29 <= R1904;
    end
    if(T2106) begin
      useRAS_28 <= R1904;
    end
    if(T2112) begin
      useRAS_27 <= R1904;
    end
    if(T2118) begin
      useRAS_26 <= R1904;
    end
    if(T2124) begin
      useRAS_25 <= R1904;
    end
    if(T2130) begin
      useRAS_24 <= R1904;
    end
    if(T2136) begin
      useRAS_23 <= R1904;
    end
    if(T2142) begin
      useRAS_22 <= R1904;
    end
    if(T2148) begin
      useRAS_21 <= R1904;
    end
    if(T2154) begin
      useRAS_20 <= R1904;
    end
    if(T2160) begin
      useRAS_19 <= R1904;
    end
    if(T2166) begin
      useRAS_18 <= R1904;
    end
    if(T2172) begin
      useRAS_17 <= R1904;
    end
    if(T2178) begin
      useRAS_16 <= R1904;
    end
    if(T2184) begin
      useRAS_15 <= R1904;
    end
    if(T2190) begin
      useRAS_14 <= R1904;
    end
    if(T2196) begin
      useRAS_13 <= R1904;
    end
    if(T2202) begin
      useRAS_12 <= R1904;
    end
    if(T2208) begin
      useRAS_11 <= R1904;
    end
    if(T2214) begin
      useRAS_10 <= R1904;
    end
    if(T2220) begin
      useRAS_9 <= R1904;
    end
    if(T2226) begin
      useRAS_8 <= R1904;
    end
    if(T2232) begin
      useRAS_7 <= R1904;
    end
    if(T2238) begin
      useRAS_6 <= R1904;
    end
    if(T2244) begin
      useRAS_5 <= R1904;
    end
    if(T2250) begin
      useRAS_4 <= R1904;
    end
    if(T2256) begin
      useRAS_3 <= R1904;
    end
    if(T2262) begin
      useRAS_2 <= R1904;
    end
    if(T2268) begin
      useRAS_1 <= R1904;
    end
    if(T2273) begin
      useRAS_0 <= R1904;
    end
    if (T2281)
      brIdx[T42] <= 1'h0;
  end
endmodule

module FlowThroughSerializer(
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_addr_beat,
    input [1:0] io_in_bits_client_xact_id,
    input [3:0] io_in_bits_manager_xact_id,
    input  io_in_bits_is_builtin_type,
    input [3:0] io_in_bits_g_type,
    input [127:0] io_in_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[1:0] io_out_bits_client_xact_id,
    output[3:0] io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[127:0] io_out_bits_data,
    output io_cnt,
    output io_done
);



  assign io_done = 1'h1;
  assign io_cnt = 1'h0;
  assign io_out_bits_data = io_in_bits_data;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_valid = io_in_valid;
  assign io_in_ready = io_out_ready;
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [11:0] io_req_bits_idx,
    input [19:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[31:0] io_resp_bits_data,
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[1:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data
);

  wire[127:0] T0;
  wire[16:0] T1;
  wire[2:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[25:0] T6;
  wire[25:0] T7;
  reg [31:0] s2_addr;
  wire[31:0] T8;
  wire[31:0] s1_addr;
  wire[31:0] T9;
  reg [11:0] s1_pgoff;
  wire[11:0] T10;
  wire T11;
  wire rdy;
  wire T12;
  wire T13;
  wire s2_miss;
  wire T14;
  wire s2_any_tag_hit;
  wire T15;
  wire T16;
  wire T17;
  wire s2_disparity_3;
  wire T18;
  reg  R19;
  wire T20;
  wire T21;
  wire T22;
  wire stall;
  wire T23;
  reg  s1_valid;
  wire T331;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  reg  R29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[7:0] T36;
  wire[7:0] T37;
  wire[7:0] T38;
  wire[5:0] T39;
  wire T40;
  reg [255:0] vb_array;
  wire[255:0] T332;
  wire[255:0] T41;
  wire[255:0] T42;
  wire[255:0] T43;
  wire[255:0] T44;
  wire[255:0] T45;
  wire[255:0] T46;
  wire[255:0] T47;
  wire[255:0] T48;
  wire[255:0] T49;
  wire[7:0] T50;
  wire[5:0] s2_idx;
  wire[1:0] repl_way;
  reg [15:0] R51;
  wire[15:0] T333;
  wire[15:0] T52;
  wire[15:0] T53;
  wire[14:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[255:0] T334;
  wire T62;
  wire[255:0] T63;
  wire[255:0] T64;
  wire T65;
  wire T66;
  reg  invalidated;
  wire T67;
  wire T68;
  wire T69;
  reg [1:0] state;
  wire[1:0] T335;
  wire[1:0] T70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire refill_done;
  wire refill_wrap;
  wire T81;
  reg [1:0] refill_cnt;
  wire[1:0] T336;
  wire[1:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire[255:0] T86;
  wire[255:0] T337;
  wire[127:0] T87;
  wire[127:0] T88;
  wire[6:0] T89;
  wire[127:0] T338;
  wire T90;
  wire[127:0] T339;
  wire T340;
  wire[255:0] T91;
  wire[255:0] T341;
  wire[127:0] T92;
  wire T93;
  wire s2_disparity_0;
  wire T94;
  reg  R95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  reg  R100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire[6:0] T107;
  wire[6:0] T108;
  wire[6:0] T109;
  wire[5:0] T110;
  wire T111;
  wire T112;
  wire[255:0] T113;
  wire[255:0] T342;
  wire[127:0] T114;
  wire[127:0] T115;
  wire[6:0] T116;
  wire[127:0] T343;
  wire T117;
  wire[127:0] T344;
  wire T345;
  wire[255:0] T118;
  wire[255:0] T346;
  wire[127:0] T119;
  wire T120;
  wire s2_disparity_1;
  wire T121;
  reg  R122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  reg  R127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[6:0] T134;
  wire[6:0] T135;
  wire[6:0] T136;
  wire[5:0] T137;
  wire T138;
  wire T139;
  wire[255:0] T140;
  wire[255:0] T141;
  wire[255:0] T142;
  wire[7:0] T143;
  wire[255:0] T347;
  wire T144;
  wire[255:0] T145;
  wire[255:0] T146;
  wire T147;
  wire s2_disparity_2;
  wire T148;
  reg  R149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  reg  R154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire[7:0] T161;
  wire[7:0] T162;
  wire[7:0] T163;
  wire[5:0] T164;
  wire T165;
  wire T166;
  wire[255:0] T167;
  wire[255:0] T168;
  wire[255:0] T169;
  wire[7:0] T170;
  wire[255:0] T348;
  wire T171;
  wire[255:0] T172;
  wire[255:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire s2_tag_hit_3;
  wire T179;
  reg  R180;
  wire T181;
  wire s1_tag_match_3;
  wire T182;
  wire[19:0] s1_tag;
  wire[19:0] T183;
  wire[79:0] T184;
  wire T207;
  wire s0_valid;
  wire T208;
  wire T209;
  wire[5:0] T205;
  wire[11:0] s0_pgoff;
  wire T206;
  wire[79:0] T185;
  wire[79:0] T186;
  wire[79:0] T187;
  wire[39:0] T188;
  wire[19:0] T189;
  wire[19:0] T349;
  wire T190;
  wire[19:0] T191;
  wire[19:0] T350;
  wire T192;
  wire[39:0] T193;
  wire[19:0] T194;
  wire[19:0] T351;
  wire T195;
  wire[19:0] T196;
  wire[19:0] T352;
  wire T197;
  wire[79:0] T198;
  wire[79:0] T199;
  wire[39:0] T200;
  wire[19:0] T201;
  wire[19:0] s2_tag;
  wire[39:0] T202;
  reg [5:0] R203;
  wire[5:0] T204;
  wire T210;
  wire s2_tag_hit_2;
  wire T211;
  reg  R212;
  wire T213;
  wire s1_tag_match_2;
  wire T214;
  wire[19:0] T215;
  wire T216;
  wire s2_tag_hit_1;
  wire T217;
  reg  R218;
  wire T219;
  wire s1_tag_match_1;
  wire T220;
  wire[19:0] T221;
  wire s2_tag_hit_0;
  wire T222;
  reg  R223;
  wire T224;
  wire s1_tag_match_0;
  wire T225;
  wire[19:0] T226;
  reg  s2_valid;
  wire T353;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire[127:0] T237;
  wire[127:0] T238;
  reg [127:0] s2_dout_3;
  wire[127:0] T239;
  wire[127:0] T240;
  wire T250;
  wire T251;
  wire T244;
  wire T245;
  wire[7:0] T249;
  wire[127:0] T242;
  wire[127:0] T243;
  wire[7:0] T246;
  reg [7:0] R247;
  wire[7:0] T248;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[127:0] T256;
  wire[127:0] T257;
  reg [127:0] s2_dout_2;
  wire[127:0] T258;
  wire[127:0] T259;
  wire T269;
  wire T270;
  wire T263;
  wire T264;
  wire[7:0] T268;
  wire[127:0] T261;
  wire[127:0] T262;
  wire[7:0] T265;
  reg [7:0] R266;
  wire[7:0] T267;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire[127:0] T275;
  wire[127:0] T276;
  reg [127:0] s2_dout_1;
  wire[127:0] T277;
  wire[127:0] T278;
  wire T288;
  wire T289;
  wire T282;
  wire T283;
  wire[7:0] T287;
  wire[127:0] T280;
  wire[127:0] T281;
  wire[7:0] T284;
  reg [7:0] R285;
  wire[7:0] T286;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire[127:0] T294;
  reg [127:0] s2_dout_0;
  wire[127:0] T295;
  wire[127:0] T296;
  wire T306;
  wire T307;
  wire T300;
  wire T301;
  wire[7:0] T305;
  wire[127:0] T298;
  wire[127:0] T299;
  wire[7:0] T302;
  reg [7:0] R303;
  wire[7:0] T304;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] s2_dout_word_3;
  wire[127:0] T314;
  wire[6:0] T315;
  wire[1:0] T316;
  wire[5:0] s2_offset;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] s2_dout_word_2;
  wire[127:0] T319;
  wire[6:0] T320;
  wire[1:0] T321;
  wire[31:0] T322;
  wire[31:0] T323;
  wire[31:0] s2_dout_word_1;
  wire[127:0] T324;
  wire[6:0] T325;
  wire[1:0] T326;
  wire[31:0] T327;
  wire[31:0] s2_dout_word_0;
  wire[127:0] T328;
  wire[6:0] T329;
  wire[1:0] T330;
  wire s2_hit;
  wire FlowThroughSerializer_io_in_ready;
  wire FlowThroughSerializer_io_out_valid;
  wire[127:0] FlowThroughSerializer_io_out_bits_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    s2_addr = {1{$random}};
    s1_pgoff = {1{$random}};
    R19 = {1{$random}};
    s1_valid = {1{$random}};
    R29 = {1{$random}};
    vb_array = {8{$random}};
    R51 = {1{$random}};
    invalidated = {1{$random}};
    state = {1{$random}};
    refill_cnt = {1{$random}};
    R95 = {1{$random}};
    R100 = {1{$random}};
    R122 = {1{$random}};
    R127 = {1{$random}};
    R149 = {1{$random}};
    R154 = {1{$random}};
    R180 = {1{$random}};
    R203 = {1{$random}};
    R212 = {1{$random}};
    R218 = {1{$random}};
    R223 = {1{$random}};
    s2_valid = {1{$random}};
    s2_dout_3 = {4{$random}};
    R247 = {1{$random}};
    s2_dout_2 = {4{$random}};
    R266 = {1{$random}};
    s2_dout_1 = {4{$random}};
    R285 = {1{$random}};
    s2_dout_0 = {4{$random}};
    R303 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_data = T0;
  assign T0 = 128'h0;
  assign io_mem_acquire_bits_union = T1;
  assign T1 = 17'h1c1;
  assign io_mem_acquire_bits_a_type = T2;
  assign T2 = 3'h1;
  assign io_mem_acquire_bits_is_builtin_type = T3;
  assign T3 = 1'h1;
  assign io_mem_acquire_bits_addr_beat = T4;
  assign T4 = 2'h0;
  assign io_mem_acquire_bits_client_xact_id = T5;
  assign T5 = 2'h0;
  assign io_mem_acquire_bits_addr_block = T6;
  assign T6 = T7;
  assign T7 = s2_addr >> 3'h6;
  assign T8 = T233 ? s1_addr : s2_addr;
  assign s1_addr = T9;
  assign T9 = {io_req_bits_ppn, s1_pgoff};
  assign T10 = T11 ? io_req_bits_idx : s1_pgoff;
  assign T11 = io_req_valid & rdy;
  assign rdy = T12;
  assign T12 = T232 & T13;
  assign T13 = s2_miss ^ 1'h1;
  assign s2_miss = s2_valid & T14;
  assign T14 = s2_any_tag_hit ^ 1'h1;
  assign s2_any_tag_hit = T15;
  assign T15 = T178 & T16;
  assign T16 = T17 ^ 1'h1;
  assign T17 = T176 | s2_disparity_3;
  assign s2_disparity_3 = T18;
  assign T18 = R29 & R19;
  assign T20 = T21 ? 1'h0 : R19;
  assign T21 = T23 & T22;
  assign T22 = stall ^ 1'h1;
  assign stall = io_resp_ready ^ 1'h1;
  assign T23 = s1_valid & rdy;
  assign T331 = reset ? 1'h0 : T24;
  assign T24 = T28 | T25;
  assign T25 = T27 & T26;
  assign T26 = io_req_bits_kill ^ 1'h1;
  assign T27 = s1_valid & stall;
  assign T28 = io_req_valid & rdy;
  assign T30 = T21 ? T31 : R29;
  assign T31 = T175 & T32;
  assign T32 = T33;
  assign T33 = T40 & T34;
  assign T34 = T35 - 1'h1;
  assign T35 = 1'h1 << T36;
  assign T36 = T37 + 8'h1;
  assign T37 = T38 - T38;
  assign T38 = {2'h3, T39};
  assign T39 = s1_pgoff[4'hb:3'h6];
  assign T40 = vb_array >> T38;
  assign T332 = reset ? 256'h0 : T41;
  assign T41 = T174 ? T167 : T42;
  assign T42 = T147 ? T140 : T43;
  assign T43 = T120 ? T113 : T44;
  assign T44 = T93 ? T86 : T45;
  assign T45 = io_invalidate ? 256'h0 : T46;
  assign T46 = T65 ? T47 : vb_array;
  assign T47 = T63 | T48;
  assign T48 = T334 & T49;
  assign T49 = 1'h1 << T50;
  assign T50 = {repl_way, s2_idx};
  assign s2_idx = s2_addr[4'hb:3'h6];
  assign repl_way = R51[1'h1:1'h0];
  assign T333 = reset ? 16'h1 : T52;
  assign T52 = s2_miss ? T53 : R51;
  assign T53 = {T55, T54};
  assign T54 = R51[4'hf:1'h1];
  assign T55 = T57 ^ T56;
  assign T56 = R51[3'h5:3'h5];
  assign T57 = T59 ^ T58;
  assign T58 = R51[2'h3:2'h3];
  assign T59 = T61 ^ T60;
  assign T60 = R51[2'h2:2'h2];
  assign T61 = R51[1'h0:1'h0];
  assign T334 = T62 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T62 = 1'h1;
  assign T63 = vb_array & T64;
  assign T64 = ~ T49;
  assign T65 = refill_done & T66;
  assign T66 = invalidated ^ 1'h1;
  assign T67 = T69 ? 1'h0 : T68;
  assign T68 = io_invalidate ? 1'h1 : invalidated;
  assign T69 = 2'h0 == state;
  assign T335 = reset ? 2'h0 : T70;
  assign T70 = T79 ? 2'h0 : T71;
  assign T71 = T77 ? 2'h3 : T72;
  assign T72 = T75 ? 2'h2 : T73;
  assign T73 = T74 ? 2'h1 : state;
  assign T74 = T69 & s2_miss;
  assign T75 = T76 & io_mem_acquire_ready;
  assign T76 = 2'h1 == state;
  assign T77 = T78 & io_mem_grant_valid;
  assign T78 = 2'h2 == state;
  assign T79 = T80 & refill_done;
  assign T80 = 2'h3 == state;
  assign refill_done = T85 & refill_wrap;
  assign refill_wrap = T84 & T81;
  assign T81 = refill_cnt == 2'h3;
  assign T336 = reset ? 2'h0 : T82;
  assign T82 = T84 ? T83 : refill_cnt;
  assign T83 = refill_cnt + 2'h1;
  assign T84 = 1'h1 & FlowThroughSerializer_io_out_valid;
  assign T85 = state == 2'h3;
  assign T86 = T91 | T337;
  assign T337 = {T339, T87};
  assign T87 = T338 & T88;
  assign T88 = 1'h1 << T89;
  assign T89 = {1'h0, s2_idx};
  assign T338 = T90 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T90 = 1'h0;
  assign T339 = T340 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T340 = T87[7'h7f:7'h7f];
  assign T91 = vb_array & T341;
  assign T341 = {128'h0, T92};
  assign T92 = ~ T88;
  assign T93 = s2_valid & s2_disparity_0;
  assign s2_disparity_0 = T94;
  assign T94 = R100 & R95;
  assign T96 = T97 ? 1'h0 : R95;
  assign T97 = T99 & T98;
  assign T98 = stall ^ 1'h1;
  assign T99 = s1_valid & rdy;
  assign T101 = T97 ? T102 : R100;
  assign T102 = T112 & T103;
  assign T103 = T104;
  assign T104 = T111 & T105;
  assign T105 = T106 - 1'h1;
  assign T106 = 1'h1 << T107;
  assign T107 = T108 + 7'h1;
  assign T108 = T109 - T109;
  assign T109 = {1'h0, T110};
  assign T110 = s1_pgoff[4'hb:3'h6];
  assign T111 = vb_array >> T109;
  assign T112 = io_invalidate ^ 1'h1;
  assign T113 = T118 | T342;
  assign T342 = {T344, T114};
  assign T114 = T343 & T115;
  assign T115 = 1'h1 << T116;
  assign T116 = {1'h1, s2_idx};
  assign T343 = T117 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T117 = 1'h0;
  assign T344 = T345 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T345 = T114[7'h7f:7'h7f];
  assign T118 = vb_array & T346;
  assign T346 = {128'h0, T119};
  assign T119 = ~ T115;
  assign T120 = s2_valid & s2_disparity_1;
  assign s2_disparity_1 = T121;
  assign T121 = R127 & R122;
  assign T123 = T124 ? 1'h0 : R122;
  assign T124 = T126 & T125;
  assign T125 = stall ^ 1'h1;
  assign T126 = s1_valid & rdy;
  assign T128 = T124 ? T129 : R127;
  assign T129 = T139 & T130;
  assign T130 = T131;
  assign T131 = T138 & T132;
  assign T132 = T133 - 1'h1;
  assign T133 = 1'h1 << T134;
  assign T134 = T135 + 7'h1;
  assign T135 = T136 - T136;
  assign T136 = {1'h1, T137};
  assign T137 = s1_pgoff[4'hb:3'h6];
  assign T138 = vb_array >> T136;
  assign T139 = io_invalidate ^ 1'h1;
  assign T140 = T145 | T141;
  assign T141 = T347 & T142;
  assign T142 = 1'h1 << T143;
  assign T143 = {2'h2, s2_idx};
  assign T347 = T144 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T144 = 1'h0;
  assign T145 = vb_array & T146;
  assign T146 = ~ T142;
  assign T147 = s2_valid & s2_disparity_2;
  assign s2_disparity_2 = T148;
  assign T148 = R154 & R149;
  assign T150 = T151 ? 1'h0 : R149;
  assign T151 = T153 & T152;
  assign T152 = stall ^ 1'h1;
  assign T153 = s1_valid & rdy;
  assign T155 = T151 ? T156 : R154;
  assign T156 = T166 & T157;
  assign T157 = T158;
  assign T158 = T165 & T159;
  assign T159 = T160 - 1'h1;
  assign T160 = 1'h1 << T161;
  assign T161 = T162 + 8'h1;
  assign T162 = T163 - T163;
  assign T163 = {2'h2, T164};
  assign T164 = s1_pgoff[4'hb:3'h6];
  assign T165 = vb_array >> T163;
  assign T166 = io_invalidate ^ 1'h1;
  assign T167 = T172 | T168;
  assign T168 = T348 & T169;
  assign T169 = 1'h1 << T170;
  assign T170 = {2'h3, s2_idx};
  assign T348 = T171 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T171 = 1'h0;
  assign T172 = vb_array & T173;
  assign T173 = ~ T169;
  assign T174 = s2_valid & s2_disparity_3;
  assign T175 = io_invalidate ^ 1'h1;
  assign T176 = T177 | s2_disparity_2;
  assign T177 = s2_disparity_0 | s2_disparity_1;
  assign T178 = T210 | s2_tag_hit_3;
  assign s2_tag_hit_3 = T179;
  assign T179 = R29 & R180;
  assign T181 = T21 ? s1_tag_match_3 : R180;
  assign s1_tag_match_3 = T182;
  assign T182 = T183 == s1_tag;
  assign s1_tag = s1_addr[5'h1f:4'hc];
  assign T183 = T184[7'h4f:6'h3c];
  assign T207 = T209 & s0_valid;
  assign s0_valid = io_req_valid | T208;
  assign T208 = s1_valid & stall;
  assign T209 = refill_done ^ 1'h1;
  assign T205 = s0_pgoff[4'hb:3'h6];
  assign s0_pgoff = T206 ? s1_pgoff : io_req_bits_idx;
  assign T206 = s1_valid & stall;
  ICache_tag_array tag_array (
    .CLK(clk),
    .RW0A(refill_done ? s2_idx : T205),
    .RW0E(T207 || refill_done),
    .RW0W(refill_done),
    .RW0I(T198),
    .RW0M(T186),
    .RW0O(T184)
  );
  assign T186 = T187;
  assign T187 = {T193, T188};
  assign T188 = {T191, T189};
  assign T189 = 20'h0 - T349;
  assign T349 = {19'h0, T190};
  assign T190 = repl_way == 2'h0;
  assign T191 = 20'h0 - T350;
  assign T350 = {19'h0, T192};
  assign T192 = repl_way == 2'h1;
  assign T193 = {T196, T194};
  assign T194 = 20'h0 - T351;
  assign T351 = {19'h0, T195};
  assign T195 = repl_way == 2'h2;
  assign T196 = 20'h0 - T352;
  assign T352 = {19'h0, T197};
  assign T197 = repl_way == 2'h3;
  assign T198 = T199;
  assign T199 = {T202, T200};
  assign T200 = {T201, T201};
  assign T201 = s2_tag;
  assign s2_tag = s2_addr[5'h1f:4'hc];
  assign T202 = {T201, T201};
  assign T204 = T207 ? T205 : R203;
  assign T210 = T216 | s2_tag_hit_2;
  assign s2_tag_hit_2 = T211;
  assign T211 = R154 & R212;
  assign T213 = T151 ? s1_tag_match_2 : R212;
  assign s1_tag_match_2 = T214;
  assign T214 = T215 == s1_tag;
  assign T215 = T184[6'h3b:6'h28];
  assign T216 = s2_tag_hit_0 | s2_tag_hit_1;
  assign s2_tag_hit_1 = T217;
  assign T217 = R127 & R218;
  assign T219 = T124 ? s1_tag_match_1 : R218;
  assign s1_tag_match_1 = T220;
  assign T220 = T221 == s1_tag;
  assign T221 = T184[6'h27:5'h14];
  assign s2_tag_hit_0 = T222;
  assign T222 = R100 & R223;
  assign T224 = T97 ? s1_tag_match_0 : R223;
  assign s1_tag_match_0 = T225;
  assign T225 = T226 == s1_tag;
  assign T226 = T184[5'h13:1'h0];
  assign T353 = reset ? 1'h0 : T227;
  assign T227 = T229 | T228;
  assign T228 = io_resp_valid & stall;
  assign T229 = T231 & T230;
  assign T230 = io_req_bits_kill ^ 1'h1;
  assign T231 = s1_valid & rdy;
  assign T232 = state == 2'h0;
  assign T233 = T235 & T234;
  assign T234 = stall ^ 1'h1;
  assign T235 = s1_valid & rdy;
  assign io_mem_acquire_valid = T236;
  assign T236 = state == 2'h1;
  assign io_resp_bits_datablock = T237;
  assign T237 = T256 | T238;
  assign T238 = s2_tag_hit_3 ? s2_dout_3 : 128'h0;
  assign T239 = T252 ? T240 : s2_dout_3;
  assign T250 = T251 & s0_valid;
  assign T251 = T244 ^ 1'h1;
  assign T244 = FlowThroughSerializer_io_out_valid & T245;
  assign T245 = repl_way == 2'h3;
  assign T249 = s0_pgoff[4'hb:3'h4];
  ICache_T241 T241 (
    .CLK(clk),
    .RW0A(T244 ? T246 : T249),
    .RW0E(T250 || T244),
    .RW0W(T244),
    .RW0I(T243),
    .RW0O(T240)
  );
  assign T243 = FlowThroughSerializer_io_out_bits_data;
  assign T246 = {s2_idx, refill_cnt};
  assign T248 = T250 ? T249 : R247;
  assign T252 = T253 & s1_tag_match_3;
  assign T253 = T255 & T254;
  assign T254 = stall ^ 1'h1;
  assign T255 = s1_valid & rdy;
  assign T256 = T275 | T257;
  assign T257 = s2_tag_hit_2 ? s2_dout_2 : 128'h0;
  assign T258 = T271 ? T259 : s2_dout_2;
  assign T269 = T270 & s0_valid;
  assign T270 = T263 ^ 1'h1;
  assign T263 = FlowThroughSerializer_io_out_valid & T264;
  assign T264 = repl_way == 2'h2;
  assign T268 = s0_pgoff[4'hb:3'h4];
  ICache_T241 T260 (
    .CLK(clk),
    .RW0A(T263 ? T265 : T268),
    .RW0E(T269 || T263),
    .RW0W(T263),
    .RW0I(T262),
    .RW0O(T259)
  );
  assign T262 = FlowThroughSerializer_io_out_bits_data;
  assign T265 = {s2_idx, refill_cnt};
  assign T267 = T269 ? T268 : R266;
  assign T271 = T272 & s1_tag_match_2;
  assign T272 = T274 & T273;
  assign T273 = stall ^ 1'h1;
  assign T274 = s1_valid & rdy;
  assign T275 = T294 | T276;
  assign T276 = s2_tag_hit_1 ? s2_dout_1 : 128'h0;
  assign T277 = T290 ? T278 : s2_dout_1;
  assign T288 = T289 & s0_valid;
  assign T289 = T282 ^ 1'h1;
  assign T282 = FlowThroughSerializer_io_out_valid & T283;
  assign T283 = repl_way == 2'h1;
  assign T287 = s0_pgoff[4'hb:3'h4];
  ICache_T241 T279 (
    .CLK(clk),
    .RW0A(T282 ? T284 : T287),
    .RW0E(T288 || T282),
    .RW0W(T282),
    .RW0I(T281),
    .RW0O(T278)
  );
  assign T281 = FlowThroughSerializer_io_out_bits_data;
  assign T284 = {s2_idx, refill_cnt};
  assign T286 = T288 ? T287 : R285;
  assign T290 = T291 & s1_tag_match_1;
  assign T291 = T293 & T292;
  assign T292 = stall ^ 1'h1;
  assign T293 = s1_valid & rdy;
  assign T294 = s2_tag_hit_0 ? s2_dout_0 : 128'h0;
  assign T295 = T308 ? T296 : s2_dout_0;
  assign T306 = T307 & s0_valid;
  assign T307 = T300 ^ 1'h1;
  assign T300 = FlowThroughSerializer_io_out_valid & T301;
  assign T301 = repl_way == 2'h0;
  assign T305 = s0_pgoff[4'hb:3'h4];
  ICache_T241 T297 (
    .CLK(clk),
    .RW0A(T300 ? T302 : T305),
    .RW0E(T306 || T300),
    .RW0W(T300),
    .RW0I(T299),
    .RW0O(T296)
  );
  assign T299 = FlowThroughSerializer_io_out_bits_data;
  assign T302 = {s2_idx, refill_cnt};
  assign T304 = T306 ? T305 : R303;
  assign T308 = T309 & s1_tag_match_0;
  assign T309 = T311 & T310;
  assign T310 = stall ^ 1'h1;
  assign T311 = s1_valid & rdy;
  assign io_resp_bits_data = T312;
  assign T312 = T317 | T313;
  assign T313 = s2_tag_hit_3 ? s2_dout_word_3 : 32'h0;
  assign s2_dout_word_3 = T314[5'h1f:1'h0];
  assign T314 = s2_dout_3 >> T315;
  assign T315 = T316 << 3'h5;
  assign T316 = s2_offset[2'h3:2'h2];
  assign s2_offset = s2_addr[3'h5:1'h0];
  assign T317 = T322 | T318;
  assign T318 = s2_tag_hit_2 ? s2_dout_word_2 : 32'h0;
  assign s2_dout_word_2 = T319[5'h1f:1'h0];
  assign T319 = s2_dout_2 >> T320;
  assign T320 = T321 << 3'h5;
  assign T321 = s2_offset[2'h3:2'h2];
  assign T322 = T327 | T323;
  assign T323 = s2_tag_hit_1 ? s2_dout_word_1 : 32'h0;
  assign s2_dout_word_1 = T324[5'h1f:1'h0];
  assign T324 = s2_dout_1 >> T325;
  assign T325 = T326 << 3'h5;
  assign T326 = s2_offset[2'h3:2'h2];
  assign T327 = s2_tag_hit_0 ? s2_dout_word_0 : 32'h0;
  assign s2_dout_word_0 = T328[5'h1f:1'h0];
  assign T328 = s2_dout_0 >> T329;
  assign T329 = T330 << 3'h5;
  assign T330 = s2_offset[2'h3:2'h2];
  assign io_resp_valid = s2_hit;
  assign s2_hit = s2_valid & s2_any_tag_hit;
  FlowThroughSerializer FlowThroughSerializer(
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_in_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_in_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_in_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_in_bits_g_type( io_mem_grant_bits_g_type ),
       .io_in_bits_data( io_mem_grant_bits_data ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       //.io_out_bits_addr_beat(  )
       //.io_out_bits_client_xact_id(  )
       //.io_out_bits_manager_xact_id(  )
       //.io_out_bits_is_builtin_type(  )
       //.io_out_bits_g_type(  )
       .io_out_bits_data( FlowThroughSerializer_io_out_bits_data )
       //.io_cnt(  )
       //.io_done(  )
  );

  always @(posedge clk) begin
    if(T233) begin
      s2_addr <= s1_addr;
    end
    if(T11) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(T21) begin
      R19 <= 1'h0;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T24;
    end
    if(T21) begin
      R29 <= T31;
    end
    if(reset) begin
      vb_array <= 256'h0;
    end else if(T174) begin
      vb_array <= T167;
    end else if(T147) begin
      vb_array <= T140;
    end else if(T120) begin
      vb_array <= T113;
    end else if(T93) begin
      vb_array <= T86;
    end else if(io_invalidate) begin
      vb_array <= 256'h0;
    end else if(T65) begin
      vb_array <= T47;
    end
    if(reset) begin
      R51 <= 16'h1;
    end else if(s2_miss) begin
      R51 <= T53;
    end
    if(T69) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T79) begin
      state <= 2'h0;
    end else if(T77) begin
      state <= 2'h3;
    end else if(T75) begin
      state <= 2'h2;
    end else if(T74) begin
      state <= 2'h1;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T84) begin
      refill_cnt <= T83;
    end
    if(T97) begin
      R95 <= 1'h0;
    end
    if(T97) begin
      R100 <= T102;
    end
    if(T124) begin
      R122 <= 1'h0;
    end
    if(T124) begin
      R127 <= T129;
    end
    if(T151) begin
      R149 <= 1'h0;
    end
    if(T151) begin
      R154 <= T156;
    end
    if(T21) begin
      R180 <= s1_tag_match_3;
    end
    if(T207) begin
      R203 <= T205;
    end
    if(T151) begin
      R212 <= s1_tag_match_2;
    end
    if(T124) begin
      R218 <= s1_tag_match_1;
    end
    if(T97) begin
      R223 <= s1_tag_match_0;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= T227;
    end
    if(T252) begin
      s2_dout_3 <= T240;
    end
    if(T250) begin
      R247 <= T249;
    end
    if(T271) begin
      s2_dout_2 <= T259;
    end
    if(T269) begin
      R266 <= T268;
    end
    if(T290) begin
      s2_dout_1 <= T278;
    end
    if(T288) begin
      R285 <= T287;
    end
    if(T308) begin
      s2_dout_0 <= T296;
    end
    if(T306) begin
      R303 <= T305;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input [7:0] io_clear_mask,
    input [33:0] io_tag,
    output io_hit,
    output[7:0] io_hits,
    output[7:0] io_valid_bits,
    input  io_write,
    input [33:0] io_write_tag,
    input [2:0] io_write_addr
);

  reg [7:0] vb_array;
  wire[7:0] T44;
  wire[7:0] T0;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[7:0] T4;
  wire[7:0] T45;
  wire T5;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[7:0] T8;
  wire[7:0] T9;
  wire[7:0] T10;
  wire[7:0] T11;
  wire[3:0] T12;
  wire[1:0] T13;
  wire hits_0;
  wire T14;
  wire[33:0] T15;
  reg [33:0] cam_tags [7:0];
  wire[33:0] T16;
  wire T17;
  wire hits_1;
  wire T18;
  wire[33:0] T19;
  wire T20;
  wire[1:0] T21;
  wire hits_2;
  wire T22;
  wire[33:0] T23;
  wire T24;
  wire hits_3;
  wire T25;
  wire[33:0] T26;
  wire T27;
  wire[3:0] T28;
  wire[1:0] T29;
  wire hits_4;
  wire T30;
  wire[33:0] T31;
  wire T32;
  wire hits_5;
  wire T33;
  wire[33:0] T34;
  wire T35;
  wire[1:0] T36;
  wire hits_6;
  wire T37;
  wire[33:0] T38;
  wire T39;
  wire hits_7;
  wire T40;
  wire[33:0] T41;
  wire T42;
  wire T43;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_valid_bits = vb_array;
  assign T44 = reset ? 8'h0 : T0;
  assign T0 = io_clear ? T8 : T1;
  assign T1 = io_write ? T2 : vb_array;
  assign T2 = T6 | T3;
  assign T3 = T45 & T4;
  assign T4 = 1'h1 << io_write_addr;
  assign T45 = T5 ? 8'hff : 8'h0;
  assign T5 = 1'h1;
  assign T6 = vb_array & T7;
  assign T7 = ~ T4;
  assign T8 = vb_array & T9;
  assign T9 = ~ io_clear_mask;
  assign io_hits = T10;
  assign T10 = T11;
  assign T11 = {T28, T12};
  assign T12 = {T21, T13};
  assign T13 = {hits_1, hits_0};
  assign hits_0 = T17 & T14;
  assign T14 = T15 == io_tag;
  assign T15 = cam_tags[3'h0];
  assign T17 = vb_array[1'h0:1'h0];
  assign hits_1 = T20 & T18;
  assign T18 = T19 == io_tag;
  assign T19 = cam_tags[3'h1];
  assign T20 = vb_array[1'h1:1'h1];
  assign T21 = {hits_3, hits_2};
  assign hits_2 = T24 & T22;
  assign T22 = T23 == io_tag;
  assign T23 = cam_tags[3'h2];
  assign T24 = vb_array[2'h2:2'h2];
  assign hits_3 = T27 & T25;
  assign T25 = T26 == io_tag;
  assign T26 = cam_tags[3'h3];
  assign T27 = vb_array[2'h3:2'h3];
  assign T28 = {T36, T29};
  assign T29 = {hits_5, hits_4};
  assign hits_4 = T32 & T30;
  assign T30 = T31 == io_tag;
  assign T31 = cam_tags[3'h4];
  assign T32 = vb_array[3'h4:3'h4];
  assign hits_5 = T35 & T33;
  assign T33 = T34 == io_tag;
  assign T34 = cam_tags[3'h5];
  assign T35 = vb_array[3'h5:3'h5];
  assign T36 = {hits_7, hits_6};
  assign hits_6 = T39 & T37;
  assign T37 = T38 == io_tag;
  assign T38 = cam_tags[3'h6];
  assign T39 = vb_array[3'h6:3'h6];
  assign hits_7 = T42 & T40;
  assign T40 = T41 == io_tag;
  assign T41 = cam_tags[3'h7];
  assign T42 = vb_array[3'h7:3'h7];
  assign io_hit = T43;
  assign T43 = io_hits != 8'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 8'h0;
    end else if(io_clear) begin
      vb_array <= T8;
    end else if(io_write) begin
      vb_array <= T2;
    end
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [27:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    input  io_req_bits_store,
    output io_resp_miss,
    output[19:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    output[7:0] io_resp_hit_idx,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate
);

  reg [2:0] r_refill_waddr;
  wire[2:0] T0;
  wire[2:0] repl_waddr;
  wire[2:0] T1;
  wire[3:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  reg [7:0] R9;
  wire[7:0] T10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[7:0] T13;
  wire[14:0] T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T498;
  wire[1:0] T499;
  wire T500;
  wire[1:0] T501;
  wire[1:0] T502;
  wire[3:0] T503;
  wire[3:0] T504;
  wire[3:0] T505;
  wire[1:0] T506;
  wire T507;
  wire T508;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire[7:0] T25;
  wire[10:0] T26;
  wire[7:0] T27;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire tlb_hit;
  wire tag_hit;
  wire[7:0] tag_hits;
  wire[7:0] T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire[7:0] w_array;
  wire[7:0] T36;
  wire[7:0] T37;
  wire[3:0] T38;
  wire[1:0] T39;
  reg  uw_array_0;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[7:0] T51;
  wire[2:0] T52;
  reg  uw_array_1;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  reg  uw_array_2;
  wire T57;
  wire T58;
  wire T59;
  reg  uw_array_3;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire[1:0] T64;
  reg  uw_array_4;
  wire T65;
  wire T66;
  wire T67;
  reg  uw_array_5;
  wire T68;
  wire T69;
  wire T70;
  wire[1:0] T71;
  reg  uw_array_6;
  wire T72;
  wire T73;
  wire T74;
  reg  uw_array_7;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[3:0] T80;
  wire[1:0] T81;
  reg  sw_array_0;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[7:0] T91;
  wire[2:0] T92;
  reg  sw_array_1;
  wire T93;
  wire T94;
  wire T95;
  wire[1:0] T96;
  reg  sw_array_2;
  wire T97;
  wire T98;
  wire T99;
  reg  sw_array_3;
  wire T100;
  wire T101;
  wire T102;
  wire[3:0] T103;
  wire[1:0] T104;
  reg  sw_array_4;
  wire T105;
  wire T106;
  wire T107;
  reg  sw_array_5;
  wire T108;
  wire T109;
  wire T110;
  wire[1:0] T111;
  reg  sw_array_6;
  wire T112;
  wire T113;
  wire T114;
  reg  sw_array_7;
  wire T115;
  wire T116;
  wire T117;
  wire priv_s;
  wire[1:0] priv;
  wire T118;
  wire T119;
  wire[7:0] T120;
  wire[7:0] T121;
  wire[3:0] T122;
  wire[1:0] T123;
  reg  dirty_array_0;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire[2:0] T128;
  reg  dirty_array_1;
  wire T129;
  wire T130;
  wire T131;
  wire[1:0] T132;
  reg  dirty_array_2;
  wire T133;
  wire T134;
  wire T135;
  reg  dirty_array_3;
  wire T136;
  wire T137;
  wire T138;
  wire[3:0] T139;
  wire[1:0] T140;
  reg  dirty_array_4;
  wire T141;
  wire T142;
  wire T143;
  reg  dirty_array_5;
  wire T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  reg  dirty_array_6;
  wire T148;
  wire T149;
  wire T150;
  reg  dirty_array_7;
  wire T151;
  wire T152;
  wire T153;
  wire vm_enabled;
  wire T154;
  wire T155;
  wire priv_uses_vm;
  wire T156;
  wire[2:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire[1:0] T161;
  wire[1:0] T162;
  wire T163;
  wire[1:0] T164;
  wire T165;
  wire[2:0] T509;
  wire[2:0] T510;
  wire[2:0] T511;
  wire[2:0] T512;
  wire[2:0] T513;
  wire[2:0] T514;
  wire[2:0] T515;
  wire T516;
  wire[7:0] T166;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire has_invalid_entry;
  wire T167;
  wire T168;
  wire tlb_miss;
  wire T169;
  wire bad_va;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire[33:0] T523;
  reg [34:0] r_refill_tag;
  wire[34:0] T175;
  wire[34:0] lookup_tag;
  wire[34:0] T176;
  wire T177;
  wire T178;
  reg [1:0] state;
  wire[1:0] T524;
  wire[1:0] T179;
  wire[1:0] T180;
  wire[1:0] T181;
  wire[1:0] T182;
  wire[1:0] T183;
  wire[1:0] T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire[33:0] T525;
  wire[7:0] T191;
  wire[7:0] T192;
  wire[7:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[7:0] T196;
  wire[7:0] T197;
  wire[3:0] T198;
  wire[1:0] T199;
  reg  valid_array_0;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[7:0] T204;
  wire[2:0] T205;
  reg  valid_array_1;
  wire T206;
  wire T207;
  wire T208;
  wire[1:0] T209;
  reg  valid_array_2;
  wire T210;
  wire T211;
  wire T212;
  reg  valid_array_3;
  wire T213;
  wire T214;
  wire T215;
  wire[3:0] T216;
  wire[1:0] T217;
  reg  valid_array_4;
  wire T218;
  wire T219;
  wire T220;
  reg  valid_array_5;
  wire T221;
  wire T222;
  wire T223;
  wire[1:0] T224;
  reg  valid_array_6;
  wire T225;
  wire T226;
  wire T227;
  reg  valid_array_7;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  reg  r_req_instruction;
  wire T233;
  reg  r_req_store;
  wire T234;
  wire[26:0] T526;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire[7:0] T240;
  wire[7:0] x_array;
  wire[7:0] T241;
  wire[7:0] T242;
  wire[3:0] T243;
  wire[1:0] T244;
  reg  ux_array_0;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire[2:0] T257;
  reg  ux_array_1;
  wire T258;
  wire T259;
  wire T260;
  wire[1:0] T261;
  reg  ux_array_2;
  wire T262;
  wire T263;
  wire T264;
  reg  ux_array_3;
  wire T265;
  wire T266;
  wire T267;
  wire[3:0] T268;
  wire[1:0] T269;
  reg  ux_array_4;
  wire T270;
  wire T271;
  wire T272;
  reg  ux_array_5;
  wire T273;
  wire T274;
  wire T275;
  wire[1:0] T276;
  reg  ux_array_6;
  wire T277;
  wire T278;
  wire T279;
  reg  ux_array_7;
  wire T280;
  wire T281;
  wire T282;
  wire[7:0] T283;
  wire[7:0] T284;
  wire[3:0] T285;
  wire[1:0] T286;
  reg  sx_array_0;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire[7:0] T296;
  wire[2:0] T297;
  reg  sx_array_1;
  wire T298;
  wire T299;
  wire T300;
  wire[1:0] T301;
  reg  sx_array_2;
  wire T302;
  wire T303;
  wire T304;
  reg  sx_array_3;
  wire T305;
  wire T306;
  wire T307;
  wire[3:0] T308;
  wire[1:0] T309;
  reg  sx_array_4;
  wire T310;
  wire T311;
  wire T312;
  reg  sx_array_5;
  wire T313;
  wire T314;
  wire T315;
  wire[1:0] T316;
  reg  sx_array_6;
  wire T317;
  wire T318;
  wire T319;
  reg  sx_array_7;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire[2:0] T327;
  wire[2:0] T328;
  wire[2:0] T329;
  wire T330;
  wire T331;
  wire[32:0] T527;
  wire[31:0] paddr;
  wire T332;
  wire[2:0] T333;
  wire[2:0] T334;
  wire[2:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[2:0] T339;
  wire[2:0] T340;
  wire[2:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[2:0] T345;
  wire[2:0] T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire addr_ok;
  wire T351;
  wire T352;
  wire[32:0] T528;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire[7:0] T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire[7:0] T379;
  wire[7:0] r_array;
  wire[7:0] T380;
  wire[7:0] T381;
  wire[3:0] T382;
  wire[1:0] T383;
  reg  ur_array_0;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire[7:0] T393;
  wire[2:0] T394;
  reg  ur_array_1;
  wire T395;
  wire T396;
  wire T397;
  wire[1:0] T398;
  reg  ur_array_2;
  wire T399;
  wire T400;
  wire T401;
  reg  ur_array_3;
  wire T402;
  wire T403;
  wire T404;
  wire[3:0] T405;
  wire[1:0] T406;
  reg  ur_array_4;
  wire T407;
  wire T408;
  wire T409;
  reg  ur_array_5;
  wire T410;
  wire T411;
  wire T412;
  wire[1:0] T413;
  reg  ur_array_6;
  wire T414;
  wire T415;
  wire T416;
  reg  ur_array_7;
  wire T417;
  wire T418;
  wire T419;
  wire[7:0] T420;
  wire[7:0] T421;
  wire[3:0] T422;
  wire[1:0] T423;
  reg  sr_array_0;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire[7:0] T431;
  wire[2:0] T432;
  reg  sr_array_1;
  wire T433;
  wire T434;
  wire T435;
  wire[1:0] T436;
  reg  sr_array_2;
  wire T437;
  wire T438;
  wire T439;
  reg  sr_array_3;
  wire T440;
  wire T441;
  wire T442;
  wire[3:0] T443;
  wire[1:0] T444;
  reg  sr_array_4;
  wire T445;
  wire T446;
  wire T447;
  reg  sr_array_5;
  wire T448;
  wire T449;
  wire T450;
  wire[1:0] T451;
  reg  sr_array_6;
  wire T452;
  wire T453;
  wire T454;
  reg  sr_array_7;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire[19:0] T463;
  wire[19:0] T464;
  wire[19:0] T465;
  wire[19:0] T466;
  wire[19:0] T467;
  reg [19:0] tag_ram [7:0];
  wire[19:0] T468;
  wire T469;
  wire[19:0] T470;
  wire[19:0] T471;
  wire[19:0] T472;
  wire T473;
  wire[19:0] T474;
  wire[19:0] T475;
  wire[19:0] T476;
  wire T477;
  wire[19:0] T478;
  wire[19:0] T479;
  wire[19:0] T480;
  wire T481;
  wire[19:0] T482;
  wire[19:0] T483;
  wire[19:0] T484;
  wire T485;
  wire[19:0] T486;
  wire[19:0] T487;
  wire[19:0] T488;
  wire T489;
  wire[19:0] T490;
  wire[19:0] T491;
  wire[19:0] T492;
  wire T493;
  wire[19:0] T494;
  wire[19:0] T495;
  wire T496;
  wire T497;
  wire[7:0] tag_cam_io_hits;
  wire[7:0] tag_cam_io_valid_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R9 = {1{$random}};
    uw_array_0 = {1{$random}};
    uw_array_1 = {1{$random}};
    uw_array_2 = {1{$random}};
    uw_array_3 = {1{$random}};
    uw_array_4 = {1{$random}};
    uw_array_5 = {1{$random}};
    uw_array_6 = {1{$random}};
    uw_array_7 = {1{$random}};
    sw_array_0 = {1{$random}};
    sw_array_1 = {1{$random}};
    sw_array_2 = {1{$random}};
    sw_array_3 = {1{$random}};
    sw_array_4 = {1{$random}};
    sw_array_5 = {1{$random}};
    sw_array_6 = {1{$random}};
    sw_array_7 = {1{$random}};
    dirty_array_0 = {1{$random}};
    dirty_array_1 = {1{$random}};
    dirty_array_2 = {1{$random}};
    dirty_array_3 = {1{$random}};
    dirty_array_4 = {1{$random}};
    dirty_array_5 = {1{$random}};
    dirty_array_6 = {1{$random}};
    dirty_array_7 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    valid_array_0 = {1{$random}};
    valid_array_1 = {1{$random}};
    valid_array_2 = {1{$random}};
    valid_array_3 = {1{$random}};
    valid_array_4 = {1{$random}};
    valid_array_5 = {1{$random}};
    valid_array_6 = {1{$random}};
    valid_array_7 = {1{$random}};
    r_req_instruction = {1{$random}};
    r_req_store = {1{$random}};
    ux_array_0 = {1{$random}};
    ux_array_1 = {1{$random}};
    ux_array_2 = {1{$random}};
    ux_array_3 = {1{$random}};
    ux_array_4 = {1{$random}};
    ux_array_5 = {1{$random}};
    ux_array_6 = {1{$random}};
    ux_array_7 = {1{$random}};
    sx_array_0 = {1{$random}};
    sx_array_1 = {1{$random}};
    sx_array_2 = {1{$random}};
    sx_array_3 = {1{$random}};
    sx_array_4 = {1{$random}};
    sx_array_5 = {1{$random}};
    sx_array_6 = {1{$random}};
    sx_array_7 = {1{$random}};
    ur_array_0 = {1{$random}};
    ur_array_1 = {1{$random}};
    ur_array_2 = {1{$random}};
    ur_array_3 = {1{$random}};
    ur_array_4 = {1{$random}};
    ur_array_5 = {1{$random}};
    ur_array_6 = {1{$random}};
    ur_array_7 = {1{$random}};
    sr_array_0 = {1{$random}};
    sr_array_1 = {1{$random}};
    sr_array_2 = {1{$random}};
    sr_array_3 = {1{$random}};
    sr_array_4 = {1{$random}};
    sr_array_5 = {1{$random}};
    sr_array_6 = {1{$random}};
    sr_array_7 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T168 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T509 : T1;
  assign T1 = T2[2'h2:1'h0];
  assign T2 = {T157, T3};
  assign T3 = T8 & T4;
  assign T4 = T5 - 1'h1;
  assign T5 = 1'h1 << T6;
  assign T6 = T7 + 3'h1;
  assign T7 = T157 - T157;
  assign T8 = R9 >> T157;
  assign T10 = T32 ? T11 : R9;
  assign T11 = T21 | T12;
  assign T12 = T20 ? 8'h0 : T13;
  assign T13 = T14[3'h7:1'h0];
  assign T14 = 8'h1 << T15;
  assign T15 = {T18, T16};
  assign T16 = T498[1'h1:1'h1];
  assign T498 = {T508, T499};
  assign T499 = {T507, T500};
  assign T500 = T501[1'h1:1'h1];
  assign T501 = T506 | T502;
  assign T502 = T503[1'h1:1'h0];
  assign T503 = T505 | T504;
  assign T504 = tag_cam_io_hits[2'h3:1'h0];
  assign T505 = tag_cam_io_hits[3'h7:3'h4];
  assign T506 = T503[2'h3:2'h2];
  assign T507 = T506 != 2'h0;
  assign T508 = T505 != 4'h0;
  assign T18 = {1'h1, T19};
  assign T19 = T498[2'h2:2'h2];
  assign T20 = T498[1'h0:1'h0];
  assign T21 = T23 & T22;
  assign T22 = ~ T13;
  assign T23 = T27 | T24;
  assign T24 = T16 ? 8'h0 : T25;
  assign T25 = T26[3'h7:1'h0];
  assign T26 = 8'h1 << T18;
  assign T27 = T29 & T28;
  assign T28 = ~ T25;
  assign T29 = T31 | T30;
  assign T30 = T19 ? 8'h0 : 8'h2;
  assign T31 = R9 & 8'hfd;
  assign T32 = io_req_valid & tlb_hit;
  assign tlb_hit = vm_enabled & tag_hit;
  assign tag_hit = tag_hits != 8'h0;
  assign tag_hits = tag_cam_io_hits & T33;
  assign T33 = T120 | T34;
  assign T34 = ~ T35;
  assign T35 = io_req_bits_store ? w_array : 8'h0;
  assign w_array = priv_s ? T78 : T36;
  assign T36 = T37;
  assign T37 = {T63, T38};
  assign T38 = {T56, T39};
  assign T39 = {uw_array_1, uw_array_0};
  assign T40 = T49 ? T41 : uw_array_0;
  assign T41 = T43 & T42;
  assign T42 = io_ptw_resp_bits_error ^ 1'h1;
  assign T43 = T45 & T44;
  assign T44 = io_ptw_resp_bits_pte_typ[1'h0:1'h0];
  assign T45 = T47 & T46;
  assign T46 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T47 = io_ptw_resp_bits_pte_v & T48;
  assign T48 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T49 = io_ptw_resp_valid & T50;
  assign T50 = T51[1'h0:1'h0];
  assign T51 = 1'h1 << T52;
  assign T52 = r_refill_waddr;
  assign T53 = T54 ? T41 : uw_array_1;
  assign T54 = io_ptw_resp_valid & T55;
  assign T55 = T51[1'h1:1'h1];
  assign T56 = {uw_array_3, uw_array_2};
  assign T57 = T58 ? T41 : uw_array_2;
  assign T58 = io_ptw_resp_valid & T59;
  assign T59 = T51[2'h2:2'h2];
  assign T60 = T61 ? T41 : uw_array_3;
  assign T61 = io_ptw_resp_valid & T62;
  assign T62 = T51[2'h3:2'h3];
  assign T63 = {T71, T64};
  assign T64 = {uw_array_5, uw_array_4};
  assign T65 = T66 ? T41 : uw_array_4;
  assign T66 = io_ptw_resp_valid & T67;
  assign T67 = T51[3'h4:3'h4];
  assign T68 = T69 ? T41 : uw_array_5;
  assign T69 = io_ptw_resp_valid & T70;
  assign T70 = T51[3'h5:3'h5];
  assign T71 = {uw_array_7, uw_array_6};
  assign T72 = T73 ? T41 : uw_array_6;
  assign T73 = io_ptw_resp_valid & T74;
  assign T74 = T51[3'h6:3'h6];
  assign T75 = T76 ? T41 : uw_array_7;
  assign T76 = io_ptw_resp_valid & T77;
  assign T77 = T51[3'h7:3'h7];
  assign T78 = T79;
  assign T79 = {T103, T80};
  assign T80 = {T96, T81};
  assign T81 = {sw_array_1, sw_array_0};
  assign T82 = T89 ? T83 : sw_array_0;
  assign T83 = T85 & T84;
  assign T84 = io_ptw_resp_bits_error ^ 1'h1;
  assign T85 = T87 & T86;
  assign T86 = io_ptw_resp_bits_pte_typ[1'h0:1'h0];
  assign T87 = io_ptw_resp_bits_pte_v & T88;
  assign T88 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T89 = io_ptw_resp_valid & T90;
  assign T90 = T91[1'h0:1'h0];
  assign T91 = 1'h1 << T92;
  assign T92 = r_refill_waddr;
  assign T93 = T94 ? T83 : sw_array_1;
  assign T94 = io_ptw_resp_valid & T95;
  assign T95 = T91[1'h1:1'h1];
  assign T96 = {sw_array_3, sw_array_2};
  assign T97 = T98 ? T83 : sw_array_2;
  assign T98 = io_ptw_resp_valid & T99;
  assign T99 = T91[2'h2:2'h2];
  assign T100 = T101 ? T83 : sw_array_3;
  assign T101 = io_ptw_resp_valid & T102;
  assign T102 = T91[2'h3:2'h3];
  assign T103 = {T111, T104};
  assign T104 = {sw_array_5, sw_array_4};
  assign T105 = T106 ? T83 : sw_array_4;
  assign T106 = io_ptw_resp_valid & T107;
  assign T107 = T91[3'h4:3'h4];
  assign T108 = T109 ? T83 : sw_array_5;
  assign T109 = io_ptw_resp_valid & T110;
  assign T110 = T91[3'h5:3'h5];
  assign T111 = {sw_array_7, sw_array_6};
  assign T112 = T113 ? T83 : sw_array_6;
  assign T113 = io_ptw_resp_valid & T114;
  assign T114 = T91[3'h6:3'h6];
  assign T115 = T116 ? T83 : sw_array_7;
  assign T116 = io_ptw_resp_valid & T117;
  assign T117 = T91[3'h7:3'h7];
  assign priv_s = priv == 2'h1;
  assign priv = T118 ? io_ptw_status_prv1 : io_ptw_status_prv;
  assign T118 = io_ptw_status_mprv & T119;
  assign T119 = io_req_bits_instruction ^ 1'h1;
  assign T120 = T121;
  assign T121 = {T139, T122};
  assign T122 = {T132, T123};
  assign T123 = {dirty_array_1, dirty_array_0};
  assign T124 = T125 ? io_ptw_resp_bits_pte_d : dirty_array_0;
  assign T125 = io_ptw_resp_valid & T126;
  assign T126 = T127[1'h0:1'h0];
  assign T127 = 1'h1 << T128;
  assign T128 = r_refill_waddr;
  assign T129 = T130 ? io_ptw_resp_bits_pte_d : dirty_array_1;
  assign T130 = io_ptw_resp_valid & T131;
  assign T131 = T127[1'h1:1'h1];
  assign T132 = {dirty_array_3, dirty_array_2};
  assign T133 = T134 ? io_ptw_resp_bits_pte_d : dirty_array_2;
  assign T134 = io_ptw_resp_valid & T135;
  assign T135 = T127[2'h2:2'h2];
  assign T136 = T137 ? io_ptw_resp_bits_pte_d : dirty_array_3;
  assign T137 = io_ptw_resp_valid & T138;
  assign T138 = T127[2'h3:2'h3];
  assign T139 = {T147, T140};
  assign T140 = {dirty_array_5, dirty_array_4};
  assign T141 = T142 ? io_ptw_resp_bits_pte_d : dirty_array_4;
  assign T142 = io_ptw_resp_valid & T143;
  assign T143 = T127[3'h4:3'h4];
  assign T144 = T145 ? io_ptw_resp_bits_pte_d : dirty_array_5;
  assign T145 = io_ptw_resp_valid & T146;
  assign T146 = T127[3'h5:3'h5];
  assign T147 = {dirty_array_7, dirty_array_6};
  assign T148 = T149 ? io_ptw_resp_bits_pte_d : dirty_array_6;
  assign T149 = io_ptw_resp_valid & T150;
  assign T150 = T127[3'h6:3'h6];
  assign T151 = T152 ? io_ptw_resp_bits_pte_d : dirty_array_7;
  assign T152 = io_ptw_resp_valid & T153;
  assign T153 = T127[3'h7:3'h7];
  assign vm_enabled = T155 & T154;
  assign T154 = io_req_bits_passthrough ^ 1'h1;
  assign T155 = T156 & priv_uses_vm;
  assign priv_uses_vm = priv <= 2'h1;
  assign T156 = io_ptw_status_vm[2'h3:2'h3];
  assign T157 = {T164, T158};
  assign T158 = T163 & T159;
  assign T159 = T160 - 1'h1;
  assign T160 = 1'h1 << T161;
  assign T161 = T162 + 2'h1;
  assign T162 = T164 - T164;
  assign T163 = R9 >> T164;
  assign T164 = {1'h1, T165};
  assign T165 = R9[1'h1:1'h1];
  assign T509 = T522 ? 1'h0 : T510;
  assign T510 = T521 ? 1'h1 : T511;
  assign T511 = T520 ? 2'h2 : T512;
  assign T512 = T519 ? 2'h3 : T513;
  assign T513 = T518 ? 3'h4 : T514;
  assign T514 = T517 ? 3'h5 : T515;
  assign T515 = T516 ? 3'h6 : 3'h7;
  assign T516 = T166[3'h6:3'h6];
  assign T166 = ~ tag_cam_io_valid_bits;
  assign T517 = T166[3'h5:3'h5];
  assign T518 = T166[3'h4:3'h4];
  assign T519 = T166[2'h3:2'h3];
  assign T520 = T166[2'h2:2'h2];
  assign T521 = T166[1'h1:1'h1];
  assign T522 = T166[1'h0:1'h0];
  assign has_invalid_entry = T167 ^ 1'h1;
  assign T167 = tag_cam_io_valid_bits == 8'hff;
  assign T168 = T174 & tlb_miss;
  assign tlb_miss = T172 & T169;
  assign T169 = bad_va ^ 1'h1;
  assign bad_va = T171 != T170;
  assign T170 = io_req_bits_vpn[5'h1a:5'h1a];
  assign T171 = io_req_bits_vpn[5'h1b:5'h1b];
  assign T172 = vm_enabled & T173;
  assign T173 = tag_hit ^ 1'h1;
  assign T174 = io_req_ready & io_req_valid;
  assign T523 = r_refill_tag[6'h21:1'h0];
  assign T175 = T168 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T176;
  assign T176 = {io_req_bits_asid, io_req_bits_vpn};
  assign T177 = T178 & io_ptw_resp_valid;
  assign T178 = state == 2'h2;
  assign T524 = reset ? 2'h0 : T179;
  assign T179 = io_ptw_resp_valid ? 2'h0 : T180;
  assign T180 = T189 ? 2'h3 : T181;
  assign T181 = T188 ? 2'h3 : T182;
  assign T182 = T187 ? 2'h2 : T183;
  assign T183 = T185 ? 2'h0 : T184;
  assign T184 = T168 ? 2'h1 : state;
  assign T185 = T186 & io_ptw_invalidate;
  assign T186 = state == 2'h1;
  assign T187 = T186 & io_ptw_req_ready;
  assign T188 = T187 & io_ptw_invalidate;
  assign T189 = T190 & io_ptw_invalidate;
  assign T190 = state == 2'h2;
  assign T525 = lookup_tag[6'h21:1'h0];
  assign T191 = io_ptw_invalidate ? 8'hff : T192;
  assign T192 = T195 | T193;
  assign T193 = tag_cam_io_hits & T194;
  assign T194 = ~ tag_hits;
  assign T195 = ~ T196;
  assign T196 = T197;
  assign T197 = {T216, T198};
  assign T198 = {T209, T199};
  assign T199 = {valid_array_1, valid_array_0};
  assign T200 = T202 ? T201 : valid_array_0;
  assign T201 = io_ptw_resp_bits_error ^ 1'h1;
  assign T202 = io_ptw_resp_valid & T203;
  assign T203 = T204[1'h0:1'h0];
  assign T204 = 1'h1 << T205;
  assign T205 = r_refill_waddr;
  assign T206 = T207 ? T201 : valid_array_1;
  assign T207 = io_ptw_resp_valid & T208;
  assign T208 = T204[1'h1:1'h1];
  assign T209 = {valid_array_3, valid_array_2};
  assign T210 = T211 ? T201 : valid_array_2;
  assign T211 = io_ptw_resp_valid & T212;
  assign T212 = T204[2'h2:2'h2];
  assign T213 = T214 ? T201 : valid_array_3;
  assign T214 = io_ptw_resp_valid & T215;
  assign T215 = T204[2'h3:2'h3];
  assign T216 = {T224, T217};
  assign T217 = {valid_array_5, valid_array_4};
  assign T218 = T219 ? T201 : valid_array_4;
  assign T219 = io_ptw_resp_valid & T220;
  assign T220 = T204[3'h4:3'h4];
  assign T221 = T222 ? T201 : valid_array_5;
  assign T222 = io_ptw_resp_valid & T223;
  assign T223 = T204[3'h5:3'h5];
  assign T224 = {valid_array_7, valid_array_6};
  assign T225 = T226 ? T201 : valid_array_6;
  assign T226 = io_ptw_resp_valid & T227;
  assign T227 = T204[3'h6:3'h6];
  assign T228 = T229 ? T201 : valid_array_7;
  assign T229 = io_ptw_resp_valid & T230;
  assign T230 = T204[3'h7:3'h7];
  assign T231 = io_ptw_invalidate | T232;
  assign T232 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits_fetch = r_req_instruction;
  assign T233 = T168 ? io_req_bits_instruction : r_req_instruction;
  assign io_ptw_req_bits_store = r_req_store;
  assign T234 = T168 ? io_req_bits_store : r_req_store;
  assign io_ptw_req_bits_prv = io_ptw_status_prv;
  assign io_ptw_req_bits_addr = T526;
  assign T526 = r_refill_tag[5'h1a:1'h0];
  assign io_ptw_req_valid = T235;
  assign T235 = state == 2'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_xcpt_if = T236;
  assign T236 = T323 | T237;
  assign T237 = tlb_hit & T238;
  assign T238 = T239 ^ 1'h1;
  assign T239 = T240 != 8'h0;
  assign T240 = x_array & tag_cam_io_hits;
  assign x_array = priv_s ? T283 : T241;
  assign T241 = T242;
  assign T242 = {T268, T243};
  assign T243 = {T261, T244};
  assign T244 = {ux_array_1, ux_array_0};
  assign T245 = T254 ? T246 : ux_array_0;
  assign T246 = T248 & T247;
  assign T247 = io_ptw_resp_bits_error ^ 1'h1;
  assign T248 = T250 & T249;
  assign T249 = io_ptw_resp_bits_pte_typ[1'h1:1'h1];
  assign T250 = T252 & T251;
  assign T251 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T252 = io_ptw_resp_bits_pte_v & T253;
  assign T253 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T254 = io_ptw_resp_valid & T255;
  assign T255 = T256[1'h0:1'h0];
  assign T256 = 1'h1 << T257;
  assign T257 = r_refill_waddr;
  assign T258 = T259 ? T246 : ux_array_1;
  assign T259 = io_ptw_resp_valid & T260;
  assign T260 = T256[1'h1:1'h1];
  assign T261 = {ux_array_3, ux_array_2};
  assign T262 = T263 ? T246 : ux_array_2;
  assign T263 = io_ptw_resp_valid & T264;
  assign T264 = T256[2'h2:2'h2];
  assign T265 = T266 ? T246 : ux_array_3;
  assign T266 = io_ptw_resp_valid & T267;
  assign T267 = T256[2'h3:2'h3];
  assign T268 = {T276, T269};
  assign T269 = {ux_array_5, ux_array_4};
  assign T270 = T271 ? T246 : ux_array_4;
  assign T271 = io_ptw_resp_valid & T272;
  assign T272 = T256[3'h4:3'h4];
  assign T273 = T274 ? T246 : ux_array_5;
  assign T274 = io_ptw_resp_valid & T275;
  assign T275 = T256[3'h5:3'h5];
  assign T276 = {ux_array_7, ux_array_6};
  assign T277 = T278 ? T246 : ux_array_6;
  assign T278 = io_ptw_resp_valid & T279;
  assign T279 = T256[3'h6:3'h6];
  assign T280 = T281 ? T246 : ux_array_7;
  assign T281 = io_ptw_resp_valid & T282;
  assign T282 = T256[3'h7:3'h7];
  assign T283 = T284;
  assign T284 = {T308, T285};
  assign T285 = {T301, T286};
  assign T286 = {sx_array_1, sx_array_0};
  assign T287 = T294 ? T288 : sx_array_0;
  assign T288 = T290 & T289;
  assign T289 = io_ptw_resp_bits_error ^ 1'h1;
  assign T290 = T292 & T291;
  assign T291 = io_ptw_resp_bits_pte_typ[1'h1:1'h1];
  assign T292 = io_ptw_resp_bits_pte_v & T293;
  assign T293 = 4'h4 <= io_ptw_resp_bits_pte_typ;
  assign T294 = io_ptw_resp_valid & T295;
  assign T295 = T296[1'h0:1'h0];
  assign T296 = 1'h1 << T297;
  assign T297 = r_refill_waddr;
  assign T298 = T299 ? T288 : sx_array_1;
  assign T299 = io_ptw_resp_valid & T300;
  assign T300 = T296[1'h1:1'h1];
  assign T301 = {sx_array_3, sx_array_2};
  assign T302 = T303 ? T288 : sx_array_2;
  assign T303 = io_ptw_resp_valid & T304;
  assign T304 = T296[2'h2:2'h2];
  assign T305 = T306 ? T288 : sx_array_3;
  assign T306 = io_ptw_resp_valid & T307;
  assign T307 = T296[2'h3:2'h3];
  assign T308 = {T316, T309};
  assign T309 = {sx_array_5, sx_array_4};
  assign T310 = T311 ? T288 : sx_array_4;
  assign T311 = io_ptw_resp_valid & T312;
  assign T312 = T296[3'h4:3'h4];
  assign T313 = T314 ? T288 : sx_array_5;
  assign T314 = io_ptw_resp_valid & T315;
  assign T315 = T296[3'h5:3'h5];
  assign T316 = {sx_array_7, sx_array_6};
  assign T317 = T318 ? T288 : sx_array_6;
  assign T318 = io_ptw_resp_valid & T319;
  assign T319 = T296[3'h6:3'h6];
  assign T320 = T321 ? T288 : sx_array_7;
  assign T321 = io_ptw_resp_valid & T322;
  assign T322 = T296[3'h7:3'h7];
  assign T323 = T324 | bad_va;
  assign T324 = T350 | T325;
  assign T325 = T326 ^ 1'h1;
  assign T326 = T327[1'h0:1'h0];
  assign T327 = T333 | T328;
  assign T328 = T330 ? T329 : 3'h0;
  assign T329 = 3'h6;
  assign T330 = T332 & T331;
  assign T331 = T527 < 33'h100000000;
  assign T527 = {1'h0, paddr};
  assign paddr = {io_resp_ppn, 12'h0};
  assign T332 = 32'h80000000 <= paddr;
  assign T333 = T339 | T334;
  assign T334 = T336 ? T335 : 3'h0;
  assign T335 = 3'h6;
  assign T336 = T338 & T337;
  assign T337 = paddr < 32'h40008200;
  assign T338 = 32'h40008000 <= paddr;
  assign T339 = T345 | T340;
  assign T340 = T342 ? T341 : 3'h0;
  assign T341 = 3'h6;
  assign T342 = T344 & T343;
  assign T343 = paddr < 32'h40008000;
  assign T344 = 32'h40000000 <= paddr;
  assign T345 = T347 ? T346 : 3'h0;
  assign T346 = 3'h7;
  assign T347 = T349 & T348;
  assign T348 = paddr < 32'h40000000;
  assign T349 = 32'h0 <= paddr;
  assign T350 = addr_ok ^ 1'h1;
  assign addr_ok = T354 | T351;
  assign T351 = T353 & T352;
  assign T352 = T528 < 33'h100000000;
  assign T528 = {1'h0, paddr};
  assign T353 = 32'h80000000 <= paddr;
  assign T354 = T358 | T355;
  assign T355 = T357 & T356;
  assign T356 = paddr < 32'h40008200;
  assign T357 = 32'h40008000 <= paddr;
  assign T358 = T362 | T359;
  assign T359 = T361 & T360;
  assign T360 = paddr < 32'h40008000;
  assign T361 = 32'h40000000 <= paddr;
  assign T362 = T364 & T363;
  assign T363 = paddr < 32'h40000000;
  assign T364 = 32'h0 <= paddr;
  assign io_resp_xcpt_st = T365;
  assign T365 = T370 | T366;
  assign T366 = tlb_hit & T367;
  assign T367 = T368 ^ 1'h1;
  assign T368 = T369 != 8'h0;
  assign T369 = w_array & tag_cam_io_hits;
  assign T370 = T371 | bad_va;
  assign T371 = T374 | T372;
  assign T372 = T373 ^ 1'h1;
  assign T373 = T327[1'h1:1'h1];
  assign T374 = addr_ok ^ 1'h1;
  assign io_resp_xcpt_ld = T375;
  assign T375 = T458 | T376;
  assign T376 = tlb_hit & T377;
  assign T377 = T378 ^ 1'h1;
  assign T378 = T379 != 8'h0;
  assign T379 = r_array & tag_cam_io_hits;
  assign r_array = priv_s ? T420 : T380;
  assign T380 = T381;
  assign T381 = {T405, T382};
  assign T382 = {T398, T383};
  assign T383 = {ur_array_1, ur_array_0};
  assign T384 = T391 ? T385 : ur_array_0;
  assign T385 = T387 & T386;
  assign T386 = io_ptw_resp_bits_error ^ 1'h1;
  assign T387 = T389 & T388;
  assign T388 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T389 = io_ptw_resp_bits_pte_v & T390;
  assign T390 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T391 = io_ptw_resp_valid & T392;
  assign T392 = T393[1'h0:1'h0];
  assign T393 = 1'h1 << T394;
  assign T394 = r_refill_waddr;
  assign T395 = T396 ? T385 : ur_array_1;
  assign T396 = io_ptw_resp_valid & T397;
  assign T397 = T393[1'h1:1'h1];
  assign T398 = {ur_array_3, ur_array_2};
  assign T399 = T400 ? T385 : ur_array_2;
  assign T400 = io_ptw_resp_valid & T401;
  assign T401 = T393[2'h2:2'h2];
  assign T402 = T403 ? T385 : ur_array_3;
  assign T403 = io_ptw_resp_valid & T404;
  assign T404 = T393[2'h3:2'h3];
  assign T405 = {T413, T406};
  assign T406 = {ur_array_5, ur_array_4};
  assign T407 = T408 ? T385 : ur_array_4;
  assign T408 = io_ptw_resp_valid & T409;
  assign T409 = T393[3'h4:3'h4];
  assign T410 = T411 ? T385 : ur_array_5;
  assign T411 = io_ptw_resp_valid & T412;
  assign T412 = T393[3'h5:3'h5];
  assign T413 = {ur_array_7, ur_array_6};
  assign T414 = T415 ? T385 : ur_array_6;
  assign T415 = io_ptw_resp_valid & T416;
  assign T416 = T393[3'h6:3'h6];
  assign T417 = T418 ? T385 : ur_array_7;
  assign T418 = io_ptw_resp_valid & T419;
  assign T419 = T393[3'h7:3'h7];
  assign T420 = T421;
  assign T421 = {T443, T422};
  assign T422 = {T436, T423};
  assign T423 = {sr_array_1, sr_array_0};
  assign T424 = T429 ? T425 : sr_array_0;
  assign T425 = T427 & T426;
  assign T426 = io_ptw_resp_bits_error ^ 1'h1;
  assign T427 = io_ptw_resp_bits_pte_v & T428;
  assign T428 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T429 = io_ptw_resp_valid & T430;
  assign T430 = T431[1'h0:1'h0];
  assign T431 = 1'h1 << T432;
  assign T432 = r_refill_waddr;
  assign T433 = T434 ? T425 : sr_array_1;
  assign T434 = io_ptw_resp_valid & T435;
  assign T435 = T431[1'h1:1'h1];
  assign T436 = {sr_array_3, sr_array_2};
  assign T437 = T438 ? T425 : sr_array_2;
  assign T438 = io_ptw_resp_valid & T439;
  assign T439 = T431[2'h2:2'h2];
  assign T440 = T441 ? T425 : sr_array_3;
  assign T441 = io_ptw_resp_valid & T442;
  assign T442 = T431[2'h3:2'h3];
  assign T443 = {T451, T444};
  assign T444 = {sr_array_5, sr_array_4};
  assign T445 = T446 ? T425 : sr_array_4;
  assign T446 = io_ptw_resp_valid & T447;
  assign T447 = T431[3'h4:3'h4];
  assign T448 = T449 ? T425 : sr_array_5;
  assign T449 = io_ptw_resp_valid & T450;
  assign T450 = T431[3'h5:3'h5];
  assign T451 = {sr_array_7, sr_array_6};
  assign T452 = T453 ? T425 : sr_array_6;
  assign T453 = io_ptw_resp_valid & T454;
  assign T454 = T431[3'h6:3'h6];
  assign T455 = T456 ? T425 : sr_array_7;
  assign T456 = io_ptw_resp_valid & T457;
  assign T457 = T431[3'h7:3'h7];
  assign T458 = T459 | bad_va;
  assign T459 = T462 | T460;
  assign T460 = T461 ^ 1'h1;
  assign T461 = T327[2'h2:2'h2];
  assign T462 = addr_ok ^ 1'h1;
  assign io_resp_ppn = T463;
  assign T463 = vm_enabled ? T465 : T464;
  assign T464 = io_req_bits_vpn[5'h13:1'h0];
  assign T465 = T470 | T466;
  assign T466 = T469 ? T467 : 20'h0;
  assign T467 = tag_ram[3'h7];
  assign T469 = tag_cam_io_hits[3'h7:3'h7];
  assign T470 = T474 | T471;
  assign T471 = T473 ? T472 : 20'h0;
  assign T472 = tag_ram[3'h6];
  assign T473 = tag_cam_io_hits[3'h6:3'h6];
  assign T474 = T478 | T475;
  assign T475 = T477 ? T476 : 20'h0;
  assign T476 = tag_ram[3'h5];
  assign T477 = tag_cam_io_hits[3'h5:3'h5];
  assign T478 = T482 | T479;
  assign T479 = T481 ? T480 : 20'h0;
  assign T480 = tag_ram[3'h4];
  assign T481 = tag_cam_io_hits[3'h4:3'h4];
  assign T482 = T486 | T483;
  assign T483 = T485 ? T484 : 20'h0;
  assign T484 = tag_ram[3'h3];
  assign T485 = tag_cam_io_hits[2'h3:2'h3];
  assign T486 = T490 | T487;
  assign T487 = T489 ? T488 : 20'h0;
  assign T488 = tag_ram[3'h2];
  assign T489 = tag_cam_io_hits[2'h2:2'h2];
  assign T490 = T494 | T491;
  assign T491 = T493 ? T492 : 20'h0;
  assign T492 = tag_ram[3'h1];
  assign T493 = tag_cam_io_hits[1'h1:1'h1];
  assign T494 = T496 ? T495 : 20'h0;
  assign T495 = tag_ram[3'h0];
  assign T496 = tag_cam_io_hits[1'h0:1'h0];
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T497;
  assign T497 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( T231 ),
       .io_clear_mask( T191 ),
       .io_tag( T525 ),
       //.io_hit(  )
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T177 ),
       .io_write_tag( T523 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T168) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T32) begin
      R9 <= T11;
    end
    if(T49) begin
      uw_array_0 <= T41;
    end
    if(T54) begin
      uw_array_1 <= T41;
    end
    if(T58) begin
      uw_array_2 <= T41;
    end
    if(T61) begin
      uw_array_3 <= T41;
    end
    if(T66) begin
      uw_array_4 <= T41;
    end
    if(T69) begin
      uw_array_5 <= T41;
    end
    if(T73) begin
      uw_array_6 <= T41;
    end
    if(T76) begin
      uw_array_7 <= T41;
    end
    if(T89) begin
      sw_array_0 <= T83;
    end
    if(T94) begin
      sw_array_1 <= T83;
    end
    if(T98) begin
      sw_array_2 <= T83;
    end
    if(T101) begin
      sw_array_3 <= T83;
    end
    if(T106) begin
      sw_array_4 <= T83;
    end
    if(T109) begin
      sw_array_5 <= T83;
    end
    if(T113) begin
      sw_array_6 <= T83;
    end
    if(T116) begin
      sw_array_7 <= T83;
    end
    if(T125) begin
      dirty_array_0 <= io_ptw_resp_bits_pte_d;
    end
    if(T130) begin
      dirty_array_1 <= io_ptw_resp_bits_pte_d;
    end
    if(T134) begin
      dirty_array_2 <= io_ptw_resp_bits_pte_d;
    end
    if(T137) begin
      dirty_array_3 <= io_ptw_resp_bits_pte_d;
    end
    if(T142) begin
      dirty_array_4 <= io_ptw_resp_bits_pte_d;
    end
    if(T145) begin
      dirty_array_5 <= io_ptw_resp_bits_pte_d;
    end
    if(T149) begin
      dirty_array_6 <= io_ptw_resp_bits_pte_d;
    end
    if(T152) begin
      dirty_array_7 <= io_ptw_resp_bits_pte_d;
    end
    if(T168) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T189) begin
      state <= 2'h3;
    end else if(T188) begin
      state <= 2'h3;
    end else if(T187) begin
      state <= 2'h2;
    end else if(T185) begin
      state <= 2'h0;
    end else if(T168) begin
      state <= 2'h1;
    end
    if(T202) begin
      valid_array_0 <= T201;
    end
    if(T207) begin
      valid_array_1 <= T201;
    end
    if(T211) begin
      valid_array_2 <= T201;
    end
    if(T214) begin
      valid_array_3 <= T201;
    end
    if(T219) begin
      valid_array_4 <= T201;
    end
    if(T222) begin
      valid_array_5 <= T201;
    end
    if(T226) begin
      valid_array_6 <= T201;
    end
    if(T229) begin
      valid_array_7 <= T201;
    end
    if(T168) begin
      r_req_instruction <= io_req_bits_instruction;
    end
    if(T168) begin
      r_req_store <= io_req_bits_store;
    end
    if(T254) begin
      ux_array_0 <= T246;
    end
    if(T259) begin
      ux_array_1 <= T246;
    end
    if(T263) begin
      ux_array_2 <= T246;
    end
    if(T266) begin
      ux_array_3 <= T246;
    end
    if(T271) begin
      ux_array_4 <= T246;
    end
    if(T274) begin
      ux_array_5 <= T246;
    end
    if(T278) begin
      ux_array_6 <= T246;
    end
    if(T281) begin
      ux_array_7 <= T246;
    end
    if(T294) begin
      sx_array_0 <= T288;
    end
    if(T299) begin
      sx_array_1 <= T288;
    end
    if(T303) begin
      sx_array_2 <= T288;
    end
    if(T306) begin
      sx_array_3 <= T288;
    end
    if(T311) begin
      sx_array_4 <= T288;
    end
    if(T314) begin
      sx_array_5 <= T288;
    end
    if(T318) begin
      sx_array_6 <= T288;
    end
    if(T321) begin
      sx_array_7 <= T288;
    end
    if(T391) begin
      ur_array_0 <= T385;
    end
    if(T396) begin
      ur_array_1 <= T385;
    end
    if(T400) begin
      ur_array_2 <= T385;
    end
    if(T403) begin
      ur_array_3 <= T385;
    end
    if(T408) begin
      ur_array_4 <= T385;
    end
    if(T411) begin
      ur_array_5 <= T385;
    end
    if(T415) begin
      ur_array_6 <= T385;
    end
    if(T418) begin
      ur_array_7 <= T385;
    end
    if(T429) begin
      sr_array_0 <= T425;
    end
    if(T434) begin
      sr_array_1 <= T425;
    end
    if(T438) begin
      sr_array_2 <= T425;
    end
    if(T441) begin
      sr_array_3 <= T425;
    end
    if(T446) begin
      sr_array_4 <= T425;
    end
    if(T449) begin
      sr_array_5 <= T425;
    end
    if(T453) begin
      sr_array_6 <= T425;
    end
    if(T456) begin
      sr_array_7 <= T425;
    end
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_pte_ppn;
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [39:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[39:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data_0,
    output io_cpu_resp_bits_mask,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output io_cpu_btb_resp_bits_mask,
    output io_cpu_btb_resp_bits_bridx,
    output[38:0] io_cpu_btb_resp_bits_target,
    output[5:0] io_cpu_btb_resp_bits_entry,
    output[6:0] io_cpu_btb_resp_bits_bht_history,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input  io_cpu_btb_update_bits_prediction_bits_mask,
    input  io_cpu_btb_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [5:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [38:0] io_cpu_btb_update_bits_pc,
    input [38:0] io_cpu_btb_update_bits_target,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isReturn,
    input [38:0] io_cpu_btb_update_bits_br_pc,
    input  io_cpu_bht_update_valid,
    input  io_cpu_bht_update_bits_prediction_valid,
    input  io_cpu_bht_update_bits_prediction_bits_taken,
    input  io_cpu_bht_update_bits_prediction_bits_mask,
    input  io_cpu_bht_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_bht_update_bits_prediction_bits_target,
    input [5:0] io_cpu_bht_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
    input [38:0] io_cpu_bht_update_bits_pc,
    input  io_cpu_bht_update_bits_taken,
    input  io_cpu_bht_update_bits_mispredict,
    input  io_cpu_ras_update_valid,
    input  io_cpu_ras_update_bits_isCall,
    input  io_cpu_ras_update_bits_isReturn,
    input [38:0] io_cpu_ras_update_bits_returnAddr,
    input  io_cpu_ras_update_bits_prediction_valid,
    input  io_cpu_ras_update_bits_prediction_bits_taken,
    input  io_cpu_ras_update_bits_prediction_bits_mask,
    input  io_cpu_ras_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_ras_update_bits_prediction_bits_target,
    input [5:0] io_cpu_ras_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
    input  io_cpu_invalidate,
    output[39:0] io_cpu_npc,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[1:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data
);

  wire[27:0] T0;
  wire[39:0] s1_pc;
  wire[39:0] T1;
  wire[39:0] T2;
  reg [39:0] s1_pc_;
  wire[39:0] T3;
  wire[39:0] T4;
  wire[39:0] npc;
  wire[39:0] T5;
  wire[39:0] predicted_npc;
  wire[39:0] ntpc;
  wire[38:0] T6;
  wire[36:0] T7;
  wire[39:0] ntpc_0;
  wire T8;
  wire T9;
  wire T10;
  wire[39:0] btbTarget;
  wire T11;
  reg [39:0] s2_pc;
  wire[39:0] T68;
  wire[39:0] T12;
  wire T13;
  wire T14;
  wire icmiss;
  wire T15;
  reg  s2_valid;
  wire T69;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire stall;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  reg  s1_same_block;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire s0_same_block;
  wire T30;
  wire[39:0] T31;
  wire[39:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[11:0] T70;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[38:0] T71;
  wire T47;
  wire T48;
  wire T49;
  wire[39:0] T50;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T51;
  wire T52;
  reg [6:0] s2_btb_resp_bits_bht_history;
  wire[6:0] T53;
  reg [5:0] s2_btb_resp_bits_entry;
  wire[5:0] T54;
  reg [38:0] s2_btb_resp_bits_target;
  wire[38:0] T55;
  reg  s2_btb_resp_bits_bridx;
  wire T56;
  reg  s2_btb_resp_bits_mask;
  wire T57;
  reg  s2_btb_resp_bits_taken;
  wire T58;
  reg  s2_btb_resp_valid;
  wire T72;
  wire T59;
  reg  s2_xcpt_if;
  wire T73;
  wire T60;
  wire T74;
  wire[1:0] T61;
  wire[1:0] T62;
  wire[1:0] T75;
  wire[31:0] T63;
  wire[127:0] fetch_data;
  wire[6:0] T64;
  wire[1:0] T65;
  wire T66;
  wire T67;
  wire btb_io_resp_valid;
  wire btb_io_resp_bits_taken;
  wire btb_io_resp_bits_mask;
  wire btb_io_resp_bits_bridx;
  wire[38:0] btb_io_resp_bits_target;
  wire[5:0] btb_io_resp_bits_entry;
  wire[6:0] btb_io_resp_bits_bht_history;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire icache_io_resp_valid;
  wire[127:0] icache_io_resp_bits_datablock;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_addr_block;
  wire[1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] icache_io_mem_acquire_bits_addr_beat;
  wire icache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] icache_io_mem_acquire_bits_a_type;
  wire[16:0] icache_io_mem_acquire_bits_union;
  wire[127:0] icache_io_mem_acquire_bits_data;
  wire icache_io_mem_grant_ready;
  wire tlb_io_resp_miss;
  wire[19:0] tlb_io_resp_ppn;
  wire tlb_io_resp_xcpt_if;
  wire tlb_io_ptw_req_valid;
  wire[26:0] tlb_io_ptw_req_bits_addr;
  wire[1:0] tlb_io_ptw_req_bits_prv;
  wire tlb_io_ptw_req_bits_store;
  wire tlb_io_ptw_req_bits_fetch;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s1_same_block = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_history = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_bridx = {1{$random}};
    s2_btb_resp_bits_mask = {1{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = s1_pc >> 4'hc;
  assign s1_pc = ~ T1;
  assign T1 = T2 | 40'h3;
  assign T2 = ~ s1_pc_;
  assign T3 = io_cpu_req_valid ? io_cpu_req_bits_pc : T4;
  assign T4 = T19 ? npc : s1_pc_;
  assign npc = T5;
  assign T5 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : ntpc;
  assign ntpc = {T8, T6};
  assign T6 = {T7, 2'h0};
  assign T7 = ntpc_0[6'h26:2'h2];
  assign ntpc_0 = s1_pc + 40'h4;
  assign T8 = T10 & T9;
  assign T9 = ntpc_0[6'h26:6'h26];
  assign T10 = s1_pc[6'h26:6'h26];
  assign btbTarget = {T11, btb_io_resp_bits_target};
  assign T11 = btb_io_resp_bits_target[6'h26:6'h26];
  assign T68 = reset ? 40'h200 : T12;
  assign T12 = T13 ? s1_pc : s2_pc;
  assign T13 = T19 & T14;
  assign T14 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T15;
  assign T15 = icache_io_resp_valid ^ 1'h1;
  assign T69 = reset ? 1'h1 : T16;
  assign T16 = io_cpu_req_valid ? 1'h0 : T17;
  assign T17 = T19 ? T18 : s2_valid;
  assign T18 = icmiss ^ 1'h1;
  assign T19 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T20;
  assign T20 = io_cpu_resp_ready ^ 1'h1;
  assign T21 = T23 & T22;
  assign T22 = icmiss ^ 1'h1;
  assign T23 = stall ^ 1'h1;
  assign T24 = T38 & T25;
  assign T25 = s1_same_block ^ 1'h1;
  assign T26 = io_cpu_req_valid ? 1'h0 : T27;
  assign T27 = T19 ? T28 : s1_same_block;
  assign T28 = s0_same_block & T29;
  assign T29 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T33 & T30;
  assign T30 = T32 == T31;
  assign T31 = s1_pc & 40'h10;
  assign T32 = ntpc & 40'h10;
  assign T33 = T35 & T34;
  assign T34 = btb_io_resp_bits_taken ^ 1'h1;
  assign T35 = T37 & T36;
  assign T36 = io_cpu_req_valid ^ 1'h1;
  assign T37 = icmiss ^ 1'h1;
  assign T38 = stall ^ 1'h1;
  assign T39 = T40 | io_ptw_invalidate;
  assign T40 = T41 | icmiss;
  assign T41 = T42 | tlb_io_resp_xcpt_if;
  assign T42 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T70 = io_cpu_npc[4'hb:1'h0];
  assign T43 = T45 & T44;
  assign T44 = s0_same_block ^ 1'h1;
  assign T45 = stall ^ 1'h1;
  assign T46 = io_cpu_invalidate | io_ptw_invalidate;
  assign T71 = s1_pc[6'h26:1'h0];
  assign T47 = T49 & T48;
  assign T48 = icmiss ^ 1'h1;
  assign T49 = stall ^ 1'h1;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_mem_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_mem_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_mem_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_mem_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_mem_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_npc = T50;
  assign T50 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T51 = T52 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T52 = T13 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign T53 = T52 ? btb_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T54 = T52 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T55 = T52 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_bridx = s2_btb_resp_bits_bridx;
  assign T56 = T52 ? btb_io_resp_bits_bridx : s2_btb_resp_bits_bridx;
  assign io_cpu_btb_resp_bits_mask = s2_btb_resp_bits_mask;
  assign T57 = T52 ? btb_io_resp_bits_mask : s2_btb_resp_bits_mask;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T58 = T52 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T72 = reset ? 1'h0 : T59;
  assign T59 = T13 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T73 = reset ? 1'h0 : T60;
  assign T60 = T13 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_mask = T74;
  assign T74 = T61[1'h0:1'h0];
  assign T61 = s2_btb_resp_valid ? T62 : 2'h3;
  assign T62 = 2'h3 & T75;
  assign T75 = {1'h0, s2_btb_resp_bits_mask};
  assign io_cpu_resp_bits_data_0 = T63;
  assign T63 = fetch_data[5'h1f:1'h0];
  assign fetch_data = icache_io_resp_bits_datablock >> T64;
  assign T64 = T65 << 3'h5;
  assign T65 = s2_pc[2'h3:2'h2];
  assign io_cpu_resp_bits_pc = s2_pc;
  assign io_cpu_resp_valid = T66;
  assign T66 = s2_valid & T67;
  assign T67 = s2_xcpt_if | icache_io_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req_valid( T47 ),
       .io_req_bits_addr( T71 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_mask( btb_io_resp_bits_mask ),
       .io_resp_bits_bridx( btb_io_resp_bits_bridx ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_history( btb_io_resp_bits_bht_history ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_btb_update_valid( io_cpu_btb_update_valid ),
       .io_btb_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_btb_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_btb_update_bits_prediction_bits_mask( io_cpu_btb_update_bits_prediction_bits_mask ),
       .io_btb_update_bits_prediction_bits_bridx( io_cpu_btb_update_bits_prediction_bits_bridx ),
       .io_btb_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_btb_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_btb_update_bits_prediction_bits_bht_history( io_cpu_btb_update_bits_prediction_bits_bht_history ),
       .io_btb_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_btb_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_btb_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_btb_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_btb_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_btb_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_btb_update_bits_br_pc( io_cpu_btb_update_bits_br_pc ),
       .io_bht_update_valid( io_cpu_bht_update_valid ),
       .io_bht_update_bits_prediction_valid( io_cpu_bht_update_bits_prediction_valid ),
       .io_bht_update_bits_prediction_bits_taken( io_cpu_bht_update_bits_prediction_bits_taken ),
       .io_bht_update_bits_prediction_bits_mask( io_cpu_bht_update_bits_prediction_bits_mask ),
       .io_bht_update_bits_prediction_bits_bridx( io_cpu_bht_update_bits_prediction_bits_bridx ),
       .io_bht_update_bits_prediction_bits_target( io_cpu_bht_update_bits_prediction_bits_target ),
       .io_bht_update_bits_prediction_bits_entry( io_cpu_bht_update_bits_prediction_bits_entry ),
       .io_bht_update_bits_prediction_bits_bht_history( io_cpu_bht_update_bits_prediction_bits_bht_history ),
       .io_bht_update_bits_prediction_bits_bht_value( io_cpu_bht_update_bits_prediction_bits_bht_value ),
       .io_bht_update_bits_pc( io_cpu_bht_update_bits_pc ),
       .io_bht_update_bits_taken( io_cpu_bht_update_bits_taken ),
       .io_bht_update_bits_mispredict( io_cpu_bht_update_bits_mispredict ),
       .io_ras_update_valid( io_cpu_ras_update_valid ),
       .io_ras_update_bits_isCall( io_cpu_ras_update_bits_isCall ),
       .io_ras_update_bits_isReturn( io_cpu_ras_update_bits_isReturn ),
       .io_ras_update_bits_returnAddr( io_cpu_ras_update_bits_returnAddr ),
       .io_ras_update_bits_prediction_valid( io_cpu_ras_update_bits_prediction_valid ),
       .io_ras_update_bits_prediction_bits_taken( io_cpu_ras_update_bits_prediction_bits_taken ),
       .io_ras_update_bits_prediction_bits_mask( io_cpu_ras_update_bits_prediction_bits_mask ),
       .io_ras_update_bits_prediction_bits_bridx( io_cpu_ras_update_bits_prediction_bits_bridx ),
       .io_ras_update_bits_prediction_bits_target( io_cpu_ras_update_bits_prediction_bits_target ),
       .io_ras_update_bits_prediction_bits_entry( io_cpu_ras_update_bits_prediction_bits_entry ),
       .io_ras_update_bits_prediction_bits_bht_history( io_cpu_ras_update_bits_prediction_bits_bht_history ),
       .io_ras_update_bits_prediction_bits_bht_value( io_cpu_ras_update_bits_prediction_bits_bht_value ),
       .io_invalidate( T46 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T43 ),
       .io_req_bits_idx( T70 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T39 ),
       .io_resp_ready( T24 ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( icache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( icache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( icache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( icache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( icache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( icache_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( icache_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T21 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T0 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_req_bits_store( 1'h0 ),
       .io_resp_miss( tlb_io_resp_miss ),
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       //.io_resp_hit_idx(  )
       .io_ptw_req_ready( io_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( tlb_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( tlb_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( tlb_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( tlb_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( io_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_ptw_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( io_ptw_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( io_ptw_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( io_ptw_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( io_ptw_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( io_ptw_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( io_ptw_resp_bits_pte_v ),
       .io_ptw_status_sd( io_ptw_status_sd ),
       .io_ptw_status_zero2( io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( io_ptw_status_zero1 ),
       .io_ptw_status_vm( io_ptw_status_vm ),
       .io_ptw_status_mprv( io_ptw_status_mprv ),
       .io_ptw_status_xs( io_ptw_status_xs ),
       .io_ptw_status_fs( io_ptw_status_fs ),
       .io_ptw_status_prv3( io_ptw_status_prv3 ),
       .io_ptw_status_ie3( io_ptw_status_ie3 ),
       .io_ptw_status_prv2( io_ptw_status_prv2 ),
       .io_ptw_status_ie2( io_ptw_status_ie2 ),
       .io_ptw_status_prv1( io_ptw_status_prv1 ),
       .io_ptw_status_ie1( io_ptw_status_ie1 ),
       .io_ptw_status_prv( io_ptw_status_prv ),
       .io_ptw_status_ie( io_ptw_status_ie ),
       .io_ptw_invalidate( io_ptw_invalidate )
  );

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T19) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 40'h200;
    end else if(T13) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T19) begin
      s2_valid <= T18;
    end
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T19) begin
      s1_same_block <= T28;
    end
    if(T52) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T52) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if(T52) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T52) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T52) begin
      s2_btb_resp_bits_bridx <= btb_io_resp_bits_bridx;
    end
    if(T52) begin
      s2_btb_resp_bits_mask <= btb_io_resp_bits_mask;
    end
    if(T52) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T13) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T13) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [1:0] io_req_bits_addr_beat,
    input [25:0] io_req_bits_addr_block,
    input [1:0] io_req_bits_client_xact_id,
    input [2:0] io_req_bits_r_type,
    input  io_req_bits_voluntary,
    input [127:0] io_req_bits_data,
    input [3:0] io_req_bits_way_en,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output[3:0] io_data_req_bits_way_en,
    output[11:0] io_data_req_bits_addr,
    input [127:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[1:0] io_release_bits_addr_beat,
    output[25:0] io_release_bits_addr_block,
    output[1:0] io_release_bits_client_xact_id,
    output[2:0] io_release_bits_r_type,
    output io_release_bits_voluntary,
    output[127:0] io_release_bits_data
);

  reg  req_voluntary;
  wire T0;
  wire T1;
  reg [2:0] req_r_type;
  wire[2:0] T2;
  reg [1:0] req_client_xact_id;
  wire[1:0] T3;
  reg [25:0] req_addr_block;
  wire[25:0] T4;
  reg [1:0] beat_cnt;
  wire[1:0] T40;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  reg  r2_data_req_fired;
  wire T41;
  wire T9;
  wire T10;
  reg  r1_data_req_fired;
  wire T42;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg  active;
  wire T43;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg [2:0] data_req_cnt;
  wire[2:0] T44;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T45;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire[11:0] T33;
  wire[7:0] T34;
  wire[1:0] T35;
  wire[5:0] req_idx;
  reg [3:0] req_way_en;
  wire[3:0] T36;
  wire fire;
  wire T37;
  wire[19:0] T38;
  wire T39;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_voluntary = {1{$random}};
    req_r_type = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr_block = {1{$random}};
    beat_cnt = {1{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    data_req_cnt = {1{$random}};
    req_way_en = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_release_bits_data = io_data_resp;
  assign io_release_bits_voluntary = req_voluntary;
  assign T0 = T1 ? io_req_bits_voluntary : req_voluntary;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_r_type = req_r_type;
  assign T2 = T1 ? io_req_bits_r_type : req_r_type;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T3 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr_block = req_addr_block;
  assign T4 = T1 ? io_req_bits_addr_block : req_addr_block;
  assign io_release_bits_addr_beat = beat_cnt;
  assign T40 = reset ? 2'h0 : T5;
  assign T5 = T7 ? T6 : beat_cnt;
  assign T6 = beat_cnt + 2'h1;
  assign T7 = io_release_ready & io_release_valid;
  assign io_release_valid = T8;
  assign T8 = active & r2_data_req_fired;
  assign T41 = reset ? 1'h0 : T9;
  assign T9 = T18 ? 1'h0 : T10;
  assign T10 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T42 = reset ? 1'h0 : T11;
  assign T11 = T18 ? 1'h0 : T12;
  assign T12 = T14 ? 1'h1 : T13;
  assign T13 = active ? 1'h0 : r1_data_req_fired;
  assign T14 = active & T15;
  assign T15 = T17 & T16;
  assign T16 = io_meta_read_ready & io_meta_read_valid;
  assign T17 = io_data_req_ready & io_data_req_valid;
  assign T18 = T8 & T19;
  assign T19 = io_release_ready ^ 1'h1;
  assign T43 = reset ? 1'h0 : T20;
  assign T20 = T1 ? 1'h1 : T21;
  assign T21 = T31 ? T22 : active;
  assign T22 = T24 | T23;
  assign T23 = io_release_ready ^ 1'h1;
  assign T24 = data_req_cnt < 3'h4;
  assign T44 = reset ? 3'h0 : T25;
  assign T25 = T1 ? 3'h0 : T26;
  assign T26 = T18 ? T29 : T27;
  assign T27 = T14 ? T28 : data_req_cnt;
  assign T28 = data_req_cnt + 3'h1;
  assign T29 = data_req_cnt - T45;
  assign T45 = {1'h0, T30};
  assign T30 = r1_data_req_fired ? 2'h2 : 2'h1;
  assign T31 = T8 & T32;
  assign T32 = r1_data_req_fired ^ 1'h1;
  assign io_data_req_bits_addr = T33;
  assign T33 = T34 << 3'h4;
  assign T34 = {req_idx, T35};
  assign T35 = data_req_cnt[1'h1:1'h0];
  assign req_idx = req_addr_block[3'h5:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T36 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T37;
  assign T37 = data_req_cnt < 3'h4;
  assign io_meta_read_bits_tag = T38;
  assign T38 = req_addr_block >> 3'h6;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T39;
  assign T39 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_voluntary <= io_req_bits_voluntary;
    end
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_addr_block <= io_req_bits_addr_block;
    end
    if(reset) begin
      beat_cnt <= 2'h0;
    end else if(T7) begin
      beat_cnt <= T6;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(T18) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T18) begin
      r1_data_req_fired <= 1'h0;
    end else if(T14) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T31) begin
      active <= T22;
    end
    if(reset) begin
      data_req_cnt <= 3'h0;
    end else if(T1) begin
      data_req_cnt <= 3'h0;
    end else if(T18) begin
      data_req_cnt <= T29;
    end else if(T14) begin
      data_req_cnt <= T28;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr_block,
    input [1:0] io_req_bits_p_type,
    //input [1:0] io_req_bits_client_xact_id
    input  io_rep_ready,
    output io_rep_valid,
    output[1:0] io_rep_bits_addr_beat,
    output[25:0] io_rep_bits_addr_block,
    output[1:0] io_rep_bits_client_xact_id,
    output[2:0] io_rep_bits_r_type,
    output io_rep_bits_voluntary,
    output[127:0] io_rep_bits_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_wb_req_bits_voluntary,
    output[127:0] io_wb_req_bits_data,
    output[3:0] io_wb_req_bits_way_en,
    input [3:0] io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_block_state_state
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  reg [3:0] way_en;
  wire[3:0] T10;
  wire T11;
  reg [3:0] state;
  wire[3:0] T68;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] T27;
  wire T28;
  wire T29;
  reg [1:0] old_coh_state;
  wire[1:0] T30;
  wire tag_matches;
  wire T31;
  wire[3:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[127:0] reply_data;
  wire reply_voluntary;
  wire[2:0] reply_r_type;
  wire[2:0] T39;
  wire[2:0] T40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] miss_coh_state;
  wire T45;
  reg [1:0] req_p_type;
  wire[1:0] T46;
  wire[2:0] T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire T51;
  wire T52;
  wire[1:0] reply_client_xact_id;
  wire[25:0] reply_addr_block;
  reg [25:0] req_addr_block;
  wire[25:0] T53;
  wire[1:0] reply_addr_beat;
  wire T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[19:0] T62;
  wire[5:0] T69;
  wire T63;
  wire[19:0] T64;
  wire[5:0] T70;
  wire T65;
  wire T66;
  wire T67;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    way_en = {1{$random}};
    state = {1{$random}};
    old_coh_state = {1{$random}};
    req_p_type = {1{$random}};
    req_addr_block = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T9 | T3;
  assign T3 = T4 ^ 1'h1;
  assign T4 = T6 | T5;
  assign T5 = 3'h2 == io_rep_bits_r_type;
  assign T6 = T8 | T7;
  assign T7 = 3'h1 == io_rep_bits_r_type;
  assign T8 = 3'h0 == io_rep_bits_r_type;
  assign T9 = io_rep_valid ^ 1'h1;
  assign io_wb_req_bits_way_en = way_en;
  assign T10 = T11 ? io_way_en : way_en;
  assign T11 = state == 4'h3;
  assign T68 = reset ? 4'h0 : T12;
  assign T12 = T38 ? 4'h0 : T13;
  assign T13 = T36 ? 4'h8 : T14;
  assign T14 = T35 ? 4'h7 : T15;
  assign T15 = T33 ? T32 : T16;
  assign T16 = T31 ? T27 : T17;
  assign T17 = T25 ? 4'h1 : T18;
  assign T18 = T11 ? 4'h4 : T19;
  assign T19 = T24 ? 4'h3 : T20;
  assign T20 = T23 ? 4'h2 : T21;
  assign T21 = T22 ? 4'h1 : state;
  assign T22 = io_req_ready & io_req_valid;
  assign T23 = io_meta_read_ready & io_meta_read_valid;
  assign T24 = state == 4'h2;
  assign T25 = T11 & T26;
  assign T26 = io_mshr_rdy ^ 1'h1;
  assign T27 = T28 ? 4'h6 : 4'h5;
  assign T28 = tag_matches & T29;
  assign T29 = 2'h3 == old_coh_state;
  assign T30 = T11 ? io_block_state_state : old_coh_state;
  assign tag_matches = way_en != 4'h0;
  assign T31 = state == 4'h4;
  assign T32 = tag_matches ? 4'h8 : 4'h0;
  assign T33 = T34 & io_rep_ready;
  assign T34 = state == 4'h5;
  assign T35 = io_wb_req_ready & io_wb_req_valid;
  assign T36 = T37 & io_wb_req_ready;
  assign T37 = state == 4'h7;
  assign T38 = io_meta_write_ready & io_meta_write_valid;
  assign io_wb_req_bits_data = reply_data;
  assign reply_data = 128'h0;
  assign io_wb_req_bits_voluntary = reply_voluntary;
  assign reply_voluntary = 1'h0;
  assign io_wb_req_bits_r_type = reply_r_type;
  assign reply_r_type = T39;
  assign T39 = T52 ? T50 : T40;
  assign T40 = T49 ? T47 : T41;
  assign T41 = T45 ? T42 : 3'h3;
  assign T42 = T43 ? 3'h2 : 3'h5;
  assign T43 = 2'h3 == T44;
  assign T44 = tag_matches ? old_coh_state : miss_coh_state;
  assign miss_coh_state = 2'h0;
  assign T45 = req_p_type == 2'h2;
  assign T46 = T22 ? io_req_bits_p_type : req_p_type;
  assign T47 = T48 ? 3'h1 : 3'h4;
  assign T48 = 2'h3 == T44;
  assign T49 = req_p_type == 2'h1;
  assign T50 = T51 ? 3'h0 : 3'h3;
  assign T51 = 2'h3 == T44;
  assign T52 = req_p_type == 2'h0;
  assign io_wb_req_bits_client_xact_id = reply_client_xact_id;
  assign reply_client_xact_id = 2'h0;
  assign io_wb_req_bits_addr_block = reply_addr_block;
  assign reply_addr_block = req_addr_block;
  assign T53 = T22 ? io_req_bits_addr_block : req_addr_block;
  assign io_wb_req_bits_addr_beat = reply_addr_beat;
  assign reply_addr_beat = 2'h0;
  assign io_wb_req_valid = T54;
  assign T54 = state == 4'h6;
  assign io_meta_write_bits_data_coh_state = T55;
  assign T55 = T56;
  assign T56 = T61 ? 2'h0 : T57;
  assign T57 = T60 ? 2'h1 : T58;
  assign T58 = T59 ? old_coh_state : old_coh_state;
  assign T59 = req_p_type == 2'h2;
  assign T60 = req_p_type == 2'h1;
  assign T61 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T62;
  assign T62 = req_addr_block >> 3'h6;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T69;
  assign T69 = req_addr_block[3'h5:1'h0];
  assign io_meta_write_valid = T63;
  assign T63 = state == 4'h8;
  assign io_meta_read_bits_tag = T64;
  assign T64 = req_addr_block >> 3'h6;
  assign io_meta_read_bits_idx = T70;
  assign T70 = req_addr_block[3'h5:1'h0];
  assign io_meta_read_valid = T65;
  assign T65 = state == 4'h1;
  assign io_rep_bits_data = reply_data;
  assign io_rep_bits_voluntary = reply_voluntary;
  assign io_rep_bits_r_type = reply_r_type;
  assign io_rep_bits_client_xact_id = reply_client_xact_id;
  assign io_rep_bits_addr_block = reply_addr_block;
  assign io_rep_bits_addr_beat = reply_addr_beat;
  assign io_rep_valid = T66;
  assign T66 = state == 4'h5;
  assign io_req_ready = T67;
  assign T67 = state == 4'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "ProbeUnit should not send releases with data");
    $finish;
  end
// synthesis translate_on
`endif
    if(T11) begin
      way_en <= io_way_en;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T38) begin
      state <= 4'h0;
    end else if(T36) begin
      state <= 4'h8;
    end else if(T35) begin
      state <= 4'h7;
    end else if(T33) begin
      state <= T32;
    end else if(T31) begin
      state <= T27;
    end else if(T25) begin
      state <= 4'h1;
    end else if(T11) begin
      state <= 4'h4;
    end else if(T24) begin
      state <= 4'h3;
    end else if(T23) begin
      state <= 4'h2;
    end else if(T22) begin
      state <= 4'h1;
    end
    if(T11) begin
      old_coh_state <= io_block_state_state;
    end
    if(T22) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(T22) begin
      req_addr_block <= io_req_bits_addr_block;
    end
  end
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [19:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [19:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[19:0] io_out_bits_tag,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[19:0] T0;
  wire T1;
  wire[5:0] T2;
  wire T3;
  wire T4;
  wire T5;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T0;
  assign T0 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T1 = chosen;
  assign io_out_bits_idx = T2;
  assign T2 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T3;
  assign T3 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T4;
  assign T4 = T5 & io_out_ready;
  assign T5 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    input [19:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input [19:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[19:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[1:0] T0;
  wire T1;
  wire[19:0] T2;
  wire[3:0] T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T0;
  assign T0 = T1 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T1 = chosen;
  assign io_out_bits_data_tag = T2;
  assign T2 = T1 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T3;
  assign T3 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T4;
  assign T4 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module LockingArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [1:0] io_in_2_bits_client_xact_id,
    input [1:0] io_in_2_bits_addr_beat,
    input  io_in_2_bits_is_builtin_type,
    input [2:0] io_in_2_bits_a_type,
    input [16:0] io_in_2_bits_union,
    input [127:0] io_in_2_bits_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[127:0] io_out_bits_data,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  reg [1:0] lockIdx;
  wire[1:0] T65;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  reg  locked;
  wire T66;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  reg [1:0] R18;
  wire[1:0] T67;
  wire[1:0] T19;
  wire[127:0] T20;
  wire[127:0] T21;
  wire T22;
  wire[1:0] T23;
  wire T24;
  wire[16:0] T25;
  wire[16:0] T26;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire[25:0] T45;
  wire[25:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R18 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid ? 2'h0 : T1;
  assign T1 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T65 = reset ? 2'h2 : T2;
  assign T2 = T7 ? T3 : lockIdx;
  assign T3 = T6 ? 2'h0 : T4;
  assign T4 = T5 ? 2'h1 : 2'h2;
  assign T5 = io_in_1_ready & io_in_1_valid;
  assign T6 = io_in_0_ready & io_in_0_valid;
  assign T7 = T9 & T8;
  assign T8 = locked ^ 1'h1;
  assign T9 = T12 & T10;
  assign T10 = io_out_bits_is_builtin_type & T11;
  assign T11 = 3'h3 == io_out_bits_a_type;
  assign T12 = io_out_ready & io_out_valid;
  assign T66 = reset ? 1'h0 : T13;
  assign T13 = T15 ? 1'h0 : T14;
  assign T14 = T7 ? 1'h1 : locked;
  assign T15 = T12 & T16;
  assign T16 = T17 == 2'h0;
  assign T17 = R18 + 2'h1;
  assign T67 = reset ? 2'h0 : T19;
  assign T19 = T9 ? T17 : R18;
  assign io_out_bits_data = T20;
  assign T20 = T24 ? io_in_2_bits_data : T21;
  assign T21 = T22 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T22 = T23[1'h0:1'h0];
  assign T23 = chosen;
  assign T24 = T23[1'h1:1'h1];
  assign io_out_bits_union = T25;
  assign T25 = T28 ? io_in_2_bits_union : T26;
  assign T26 = T27 ? io_in_1_bits_union : io_in_0_bits_union;
  assign T27 = T23[1'h0:1'h0];
  assign T28 = T23[1'h1:1'h1];
  assign io_out_bits_a_type = T29;
  assign T29 = T32 ? io_in_2_bits_a_type : T30;
  assign T30 = T31 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign T31 = T23[1'h0:1'h0];
  assign T32 = T23[1'h1:1'h1];
  assign io_out_bits_is_builtin_type = T33;
  assign T33 = T36 ? io_in_2_bits_is_builtin_type : T34;
  assign T34 = T35 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T35 = T23[1'h0:1'h0];
  assign T36 = T23[1'h1:1'h1];
  assign io_out_bits_addr_beat = T37;
  assign T37 = T40 ? io_in_2_bits_addr_beat : T38;
  assign T38 = T39 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T39 = T23[1'h0:1'h0];
  assign T40 = T23[1'h1:1'h1];
  assign io_out_bits_client_xact_id = T41;
  assign T41 = T44 ? io_in_2_bits_client_xact_id : T42;
  assign T42 = T43 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T43 = T23[1'h0:1'h0];
  assign T44 = T23[1'h1:1'h1];
  assign io_out_bits_addr_block = T45;
  assign T45 = T48 ? io_in_2_bits_addr_block : T46;
  assign T46 = T47 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T47 = T23[1'h0:1'h0];
  assign T48 = T23[1'h1:1'h1];
  assign io_out_valid = T49;
  assign T49 = T52 ? io_in_2_valid : T50;
  assign T50 = T51 ? io_in_1_valid : io_in_0_valid;
  assign T51 = T23[1'h0:1'h0];
  assign T52 = T23[1'h1:1'h1];
  assign io_in_0_ready = T53;
  assign T53 = T54 & io_out_ready;
  assign T54 = locked ? T55 : 1'h1;
  assign T55 = lockIdx == 2'h0;
  assign io_in_1_ready = T56;
  assign T56 = T57 & io_out_ready;
  assign T57 = locked ? T59 : T58;
  assign T58 = io_in_0_valid ^ 1'h1;
  assign T59 = lockIdx == 2'h1;
  assign io_in_2_ready = T60;
  assign T60 = T61 & io_out_ready;
  assign T61 = locked ? T64 : T62;
  assign T62 = T63 ^ 1'h1;
  assign T63 = io_in_0_valid | io_in_1_valid;
  assign T64 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T7) begin
      lockIdx <= T3;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h0;
    end else if(T7) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T9) begin
      R18 <= T17;
    end
  end
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_r_type,
    input  io_in_1_bits_voluntary,
    input [127:0] io_in_1_bits_data,
    input [3:0] io_in_1_bits_way_en,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_r_type,
    input  io_in_0_bits_voluntary,
    input [127:0] io_in_0_bits_data,
    input [3:0] io_in_0_bits_way_en,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_r_type,
    output io_out_bits_voluntary,
    output[127:0] io_out_bits_data,
    output[3:0] io_out_bits_way_en,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[3:0] T0;
  wire T1;
  wire[127:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[1:0] T5;
  wire[25:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_way_en = T0;
  assign T0 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T1 = chosen;
  assign io_out_bits_data = T2;
  assign T2 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_voluntary = T3;
  assign T3 = T1 ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign io_out_bits_r_type = T4;
  assign T4 = T1 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign io_out_bits_client_xact_id = T5;
  assign T5 = T1 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T6;
  assign T6 = T1 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_bits_addr_beat = T7;
  assign T7 = T1 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_7(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [39:0] io_in_1_bits_addr,
    input [8:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_kill,
    input  io_in_1_bits_phys,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [39:0] io_in_0_bits_addr,
    input [8:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_kill,
    input  io_in_0_bits_phys,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output[39:0] io_out_bits_addr,
    output[8:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[2:0] io_out_bits_typ,
    output io_out_bits_kill,
    output io_out_bits_phys,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[4:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] T4;
  wire[4:0] T5;
  wire[8:0] T6;
  wire[39:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T0;
  assign T0 = T1 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T1 = chosen;
  assign io_out_bits_phys = T2;
  assign T2 = T1 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_kill = T3;
  assign T3 = T1 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_bits_typ = T4;
  assign T4 = T1 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_cmd = T5;
  assign T5 = T1 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T6;
  assign T6 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_addr = T7;
  assign T7 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_8(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits = T0;
  assign T0 = T1 ? io_in_1_bits : io_in_0_bits;
  assign T1 = chosen;
  assign io_out_valid = T2;
  assign T2 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T3;
  assign T3 = T4 & io_out_ready;
  assign T4 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_14(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [39:0] io_enq_bits_addr,
    input [8:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_kill,
    input  io_enq_bits_phys,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[39:0] io_deq_bits_addr,
    output[8:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_kill,
    output io_deq_bits_phys,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T29;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  reg [3:0] R4;
  wire[3:0] T30;
  wire[3:0] T5;
  wire[3:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T31;
  wire T8;
  wire T9;
  wire[4:0] T10;
  wire[63:0] T11;
  reg [63:0] ram [15:0];
  wire[63:0] T12;
  wire[63:0] T13;
  wire[63:0] T14;
  wire[9:0] T15;
  wire[5:0] T16;
  wire[3:0] T17;
  wire[53:0] T18;
  wire[13:0] T19;
  wire T20;
  wire T21;
  wire[2:0] T22;
  wire[4:0] T23;
  wire[8:0] T24;
  wire[39:0] T25;
  wire T26;
  wire empty;
  wire T27;
  wire T28;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T29 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T30 = reset ? 4'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T31 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T10;
  assign T10 = T11[3'h4:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_phys, io_enq_bits_sdq_id};
  assign T17 = {io_enq_bits_typ, io_enq_bits_kill};
  assign T18 = {io_enq_bits_addr, T19};
  assign T19 = {io_enq_bits_tag, io_enq_bits_cmd};
  assign io_deq_bits_phys = T20;
  assign T20 = T11[3'h5:3'h5];
  assign io_deq_bits_kill = T21;
  assign T21 = T11[3'h6:3'h6];
  assign io_deq_bits_typ = T22;
  assign T22 = T11[4'h9:3'h7];
  assign io_deq_bits_cmd = T23;
  assign T23 = T11[4'he:4'ha];
  assign io_deq_bits_tag = T24;
  assign T24 = T11[5'h17:4'hf];
  assign io_deq_bits_addr = T25;
  assign T25 = T11[6'h3f:5'h18];
  assign io_deq_valid = T26;
  assign T26 = empty ^ 1'h1;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 4'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input [39:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output[127:0] io_mem_req_bits_data,
    output[3:0] io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[8:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_wb_req_bits_voluntary,
    output[127:0] io_wb_req_bits_data,
    output[3:0] io_wb_req_bits_way_en,
    output io_probe_rdy
);

  wire T0;
  wire T1;
  wire T2;
  reg [3:0] state;
  wire[3:0] T216;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  wire refill_count_done;
  wire T22;
  reg [1:0] refill_cnt;
  wire[1:0] T217;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire gnt_multi_data;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire sec_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire cmd_requires_second_acquire;
  wire T80;
  wire T81;
  wire T82;
  reg [4:0] req_cmd;
  wire[4:0] T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire idx_match;
  wire[5:0] T115;
  wire[5:0] req_idx;
  reg [39:0] req_addr;
  wire[39:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg [1:0] meta_hazard;
  wire[1:0] T218;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg [3:0] req_way_en;
  wire[3:0] T133;
  wire[127:0] T134;
  wire T135;
  wire[2:0] T136;
  wire[2:0] T137;
  wire T138;
  reg [1:0] req_old_meta_coh_state;
  wire[1:0] T139;
  wire[1:0] T140;
  wire[25:0] T141;
  wire[25:0] T142;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T143;
  wire[1:0] T144;
  wire T145;
  wire[4:0] T146;
  wire[39:0] T219;
  wire[31:0] T147;
  wire[31:0] T148;
  wire[11:0] T149;
  wire[5:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  reg [1:0] new_coh_state_state;
  wire[1:0] T154;
  wire[1:0] T220;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[1:0] coh_on_grant_state;
  wire[1:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[1:0] coh_on_hit_state;
  wire[1:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[11:0] T187;
  wire[7:0] T188;
  wire[127:0] T189;
  wire[16:0] T190;
  wire[16:0] T221;
  wire[5:0] T191;
  wire[2:0] T192;
  wire[2:0] T222;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire[1:0] T205;
  wire[1:0] T206;
  wire[25:0] T207;
  wire[25:0] T208;
  wire[25:0] T209;
  wire T210;
  wire[19:0] T223;
  wire[27:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire[39:0] rpq_io_deq_bits_addr;
  wire[8:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire[4:0] rpq_io_deq_bits_sdq_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_cmd = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_coh_state = {1{$random}};
    req_old_meta_tag = {1{$random}};
    new_coh_state_state = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T69 ? 1'h0 : T1;
  assign T1 = T67 | T2;
  assign T2 = state == 4'h0;
  assign T216 = reset ? 4'h0 : T3;
  assign T3 = T65 ? T63 : T4;
  assign T4 = T61 ? 4'h4 : T5;
  assign T5 = T38 ? 4'h6 : T6;
  assign T6 = T37 ? 4'h2 : T7;
  assign T7 = T35 ? 4'h3 : T8;
  assign T8 = T33 ? 4'h4 : T9;
  assign T9 = T32 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T31 & refill_done;
  assign refill_done = io_mem_grant_valid & T21;
  assign T21 = T30 | refill_count_done;
  assign refill_count_done = T25 & T22;
  assign T22 = refill_cnt == 2'h3;
  assign T217 = reset ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_cnt;
  assign T24 = refill_cnt + 2'h1;
  assign T25 = io_mem_grant_valid & gnt_multi_data;
  assign gnt_multi_data = io_mem_grant_bits_is_builtin_type ? T29 : T26;
  assign T26 = T28 | T27;
  assign T27 = 4'h1 == io_mem_grant_bits_g_type;
  assign T28 = 4'h0 == io_mem_grant_bits_g_type;
  assign T29 = 4'h5 == io_mem_grant_bits_g_type;
  assign T30 = gnt_multi_data ^ 1'h1;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & io_mem_grant_valid;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T59 & T39;
  assign T39 = T48 ? T45 : T40;
  assign T40 = T42 | T41;
  assign T41 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T42 = T44 | T43;
  assign T43 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T44 = 2'h1 == io_req_bits_old_meta_coh_state;
  assign T45 = T47 | T46;
  assign T46 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T47 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T60 & io_req_bits_tag_match;
  assign T60 = io_req_pri_val & io_req_pri_rdy;
  assign T61 = T59 & T62;
  assign T62 = T39 ^ 1'h1;
  assign T63 = T64 ? 4'h1 : 4'h3;
  assign T64 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T65 = T60 & T66;
  assign T66 = io_req_bits_tag_match ^ 1'h1;
  assign T67 = io_replay_ready & T68;
  assign T68 = state == 4'h8;
  assign T69 = io_meta_read_ready ^ 1'h1;
  assign T70 = T75 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T74 | T73;
  assign T73 = io_req_bits_cmd == 5'h3;
  assign T74 = io_req_bits_cmd == 5'h2;
  assign T75 = T117 | T76;
  assign T76 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T77;
  assign T77 = T110 | T78;
  assign T78 = T107 & T79;
  assign T79 = cmd_requires_second_acquire ^ 1'h1;
  assign cmd_requires_second_acquire = T96 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T87 | T82;
  assign T82 = req_cmd == 5'h6;
  assign T83 = T60 ? io_req_bits_cmd : T84;
  assign T84 = T85 ? io_req_bits_cmd : req_cmd;
  assign T85 = T86 & cmd_requires_second_acquire;
  assign T86 = io_req_sec_val & io_req_sec_rdy;
  assign T87 = T89 | T88;
  assign T88 = req_cmd == 5'h3;
  assign T89 = T93 | T90;
  assign T90 = T92 | T91;
  assign T91 = req_cmd == 5'h4;
  assign T92 = req_cmd[2'h3:2'h3];
  assign T93 = T95 | T94;
  assign T94 = req_cmd == 5'h7;
  assign T95 = req_cmd == 5'h1;
  assign T96 = T98 | T97;
  assign T97 = io_req_bits_cmd == 5'h6;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h3;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3:2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign T107 = T109 | T108;
  assign T108 = 4'h5 == state;
  assign T109 = 4'h4 == state;
  assign T110 = T112 | T111;
  assign T111 = 4'h3 == state;
  assign T112 = T114 | T113;
  assign T113 = 4'h2 == state;
  assign T114 = 4'h1 == state;
  assign idx_match = req_idx == T115;
  assign T115 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T116 = T60 ? io_req_bits_addr : req_addr;
  assign T117 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T118;
  assign T118 = T132 | T119;
  assign T119 = T126 & T120;
  assign T120 = meta_hazard == 2'h0;
  assign T218 = reset ? 2'h0 : T121;
  assign T121 = T125 ? 2'h1 : T122;
  assign T122 = T124 ? T123 : meta_hazard;
  assign T123 = meta_hazard + 2'h1;
  assign T124 = meta_hazard != 2'h0;
  assign T125 = io_meta_write_ready & io_meta_write_valid;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T129 | T128;
  assign T128 = 4'h3 == state;
  assign T129 = T131 | T130;
  assign T130 = 4'h2 == state;
  assign T131 = 4'h1 == state;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T60 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_data = T134;
  assign T134 = 128'h0;
  assign io_wb_req_bits_voluntary = T135;
  assign T135 = 1'h1;
  assign io_wb_req_bits_r_type = T136;
  assign T136 = T137;
  assign T137 = T138 ? 3'h0 : 3'h3;
  assign T138 = 2'h3 == req_old_meta_coh_state;
  assign T139 = T60 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign io_wb_req_bits_client_xact_id = T140;
  assign T140 = 2'h0;
  assign io_wb_req_bits_addr_block = T141;
  assign T141 = T142;
  assign T142 = {req_old_meta_tag, req_idx};
  assign T143 = T60 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_bits_addr_beat = T144;
  assign T144 = 2'h0;
  assign io_wb_req_valid = T145;
  assign T145 = state == 4'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_cmd = T146;
  assign T146 = T69 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T219;
  assign T219 = {8'h0, T147};
  assign T147 = T148;
  assign T148 = {io_tag, T149};
  assign T149 = {req_idx, T150};
  assign T150 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_valid = T151;
  assign T151 = T152 & rpq_io_deq_valid;
  assign T152 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T153;
  assign T153 = T182 ? T181 : new_coh_state_state;
  assign T154 = 2'h0;
  assign T220 = reset ? T154 : T155;
  assign T155 = T38 ? coh_on_hit_state : T156;
  assign T156 = T172 ? coh_on_grant_state : new_coh_state_state;
  assign coh_on_grant_state = T157;
  assign T157 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T158;
  assign T158 = T171 ? 2'h1 : T159;
  assign T159 = T170 ? T162 : T160;
  assign T160 = T161 ? 2'h3 : 2'h0;
  assign T161 = io_mem_grant_bits_g_type == 4'h2;
  assign T162 = T163 ? 2'h3 : 2'h2;
  assign T163 = T167 | T164;
  assign T164 = T166 | T165;
  assign T165 = req_cmd == 5'h4;
  assign T166 = req_cmd[2'h3:2'h3];
  assign T167 = T169 | T168;
  assign T168 = req_cmd == 5'h7;
  assign T169 = req_cmd == 5'h1;
  assign T170 = io_mem_grant_bits_g_type == 4'h1;
  assign T171 = io_mem_grant_bits_g_type == 4'h0;
  assign T172 = T31 & io_mem_grant_valid;
  assign coh_on_hit_state = T173;
  assign T173 = T174 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T174 = T178 | T175;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h4;
  assign T177 = io_req_bits_cmd[2'h3:2'h3];
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h7;
  assign T180 = io_req_bits_cmd == 5'h1;
  assign T181 = 2'h0;
  assign T182 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T183;
  assign T183 = T185 | T184;
  assign T184 = state == 4'h3;
  assign T185 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T186;
  assign T186 = state == 4'h8;
  assign io_refill_addr = T187;
  assign T187 = T188 << 3'h4;
  assign T188 = {req_idx, refill_cnt};
  assign io_refill_way_en = req_way_en;
  assign io_mem_req_bits_data = T189;
  assign T189 = 128'h0;
  assign io_mem_req_bits_union = T190;
  assign T190 = T221;
  assign T221 = {11'h0, T191};
  assign T191 = {req_cmd, 1'h1};
  assign io_mem_req_bits_a_type = T192;
  assign T192 = T222;
  assign T222 = {2'h0, T193};
  assign T193 = T195 | T194;
  assign T194 = req_cmd == 5'h6;
  assign T195 = T197 | T196;
  assign T196 = req_cmd == 5'h3;
  assign T197 = T201 | T198;
  assign T198 = T200 | T199;
  assign T199 = req_cmd == 5'h4;
  assign T200 = req_cmd[2'h3:2'h3];
  assign T201 = T203 | T202;
  assign T202 = req_cmd == 5'h7;
  assign T203 = req_cmd == 5'h1;
  assign io_mem_req_bits_is_builtin_type = T204;
  assign T204 = 1'h0;
  assign io_mem_req_bits_addr_beat = T205;
  assign T205 = 2'h0;
  assign io_mem_req_bits_client_xact_id = T206;
  assign T206 = 2'h0;
  assign io_mem_req_bits_addr_block = T207;
  assign T207 = T208;
  assign T208 = T209;
  assign T209 = {io_tag, req_idx};
  assign io_mem_req_valid = T210;
  assign T210 = state == 4'h4;
  assign io_tag = T223;
  assign T223 = T211[5'h13:1'h0];
  assign T211 = req_addr >> 4'hc;
  assign io_idx_match = T212;
  assign T212 = T213 & idx_match;
  assign T213 = state != 4'h0;
  assign io_req_sec_rdy = T214;
  assign T214 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T215;
  assign T215 = state == 4'h0;
  Queue_14 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T70 ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T65) begin
      state <= T63;
    end else if(T61) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T24;
    end
    if(T60) begin
      req_cmd <= io_req_bits_cmd;
    end else if(T85) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T60) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T125) begin
      meta_hazard <= 2'h1;
    end else if(T124) begin
      meta_hazard <= T123;
    end
    if(T60) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T60) begin
      req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
    end
    if(T60) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(reset) begin
      new_coh_state_state <= T154;
    end else if(T38) begin
      new_coh_state_state <= coh_on_hit_state;
    end else if(T172) begin
      new_coh_state_state <= coh_on_grant_state;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input [39:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output[127:0] io_mem_req_bits_data,
    output[3:0] io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[8:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_wb_req_bits_voluntary,
    output[127:0] io_wb_req_bits_data,
    output[3:0] io_wb_req_bits_way_en,
    output io_probe_rdy
);

  wire T0;
  wire T1;
  wire T2;
  reg [3:0] state;
  wire[3:0] T216;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  wire refill_count_done;
  wire T22;
  reg [1:0] refill_cnt;
  wire[1:0] T217;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire gnt_multi_data;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire sec_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire cmd_requires_second_acquire;
  wire T80;
  wire T81;
  wire T82;
  reg [4:0] req_cmd;
  wire[4:0] T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire idx_match;
  wire[5:0] T115;
  wire[5:0] req_idx;
  reg [39:0] req_addr;
  wire[39:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg [1:0] meta_hazard;
  wire[1:0] T218;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg [3:0] req_way_en;
  wire[3:0] T133;
  wire[127:0] T134;
  wire T135;
  wire[2:0] T136;
  wire[2:0] T137;
  wire T138;
  reg [1:0] req_old_meta_coh_state;
  wire[1:0] T139;
  wire[1:0] T140;
  wire[25:0] T141;
  wire[25:0] T142;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T143;
  wire[1:0] T144;
  wire T145;
  wire[4:0] T146;
  wire[39:0] T219;
  wire[31:0] T147;
  wire[31:0] T148;
  wire[11:0] T149;
  wire[5:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  reg [1:0] new_coh_state_state;
  wire[1:0] T154;
  wire[1:0] T220;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[1:0] coh_on_grant_state;
  wire[1:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[1:0] coh_on_hit_state;
  wire[1:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[11:0] T187;
  wire[7:0] T188;
  wire[127:0] T189;
  wire[16:0] T190;
  wire[16:0] T221;
  wire[5:0] T191;
  wire[2:0] T192;
  wire[2:0] T222;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire[1:0] T205;
  wire[1:0] T206;
  wire[25:0] T207;
  wire[25:0] T208;
  wire[25:0] T209;
  wire T210;
  wire[19:0] T223;
  wire[27:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire[39:0] rpq_io_deq_bits_addr;
  wire[8:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire[4:0] rpq_io_deq_bits_sdq_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_cmd = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_coh_state = {1{$random}};
    req_old_meta_tag = {1{$random}};
    new_coh_state_state = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T69 ? 1'h0 : T1;
  assign T1 = T67 | T2;
  assign T2 = state == 4'h0;
  assign T216 = reset ? 4'h0 : T3;
  assign T3 = T65 ? T63 : T4;
  assign T4 = T61 ? 4'h4 : T5;
  assign T5 = T38 ? 4'h6 : T6;
  assign T6 = T37 ? 4'h2 : T7;
  assign T7 = T35 ? 4'h3 : T8;
  assign T8 = T33 ? 4'h4 : T9;
  assign T9 = T32 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T31 & refill_done;
  assign refill_done = io_mem_grant_valid & T21;
  assign T21 = T30 | refill_count_done;
  assign refill_count_done = T25 & T22;
  assign T22 = refill_cnt == 2'h3;
  assign T217 = reset ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_cnt;
  assign T24 = refill_cnt + 2'h1;
  assign T25 = io_mem_grant_valid & gnt_multi_data;
  assign gnt_multi_data = io_mem_grant_bits_is_builtin_type ? T29 : T26;
  assign T26 = T28 | T27;
  assign T27 = 4'h1 == io_mem_grant_bits_g_type;
  assign T28 = 4'h0 == io_mem_grant_bits_g_type;
  assign T29 = 4'h5 == io_mem_grant_bits_g_type;
  assign T30 = gnt_multi_data ^ 1'h1;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & io_mem_grant_valid;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T59 & T39;
  assign T39 = T48 ? T45 : T40;
  assign T40 = T42 | T41;
  assign T41 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T42 = T44 | T43;
  assign T43 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T44 = 2'h1 == io_req_bits_old_meta_coh_state;
  assign T45 = T47 | T46;
  assign T46 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T47 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T60 & io_req_bits_tag_match;
  assign T60 = io_req_pri_val & io_req_pri_rdy;
  assign T61 = T59 & T62;
  assign T62 = T39 ^ 1'h1;
  assign T63 = T64 ? 4'h1 : 4'h3;
  assign T64 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T65 = T60 & T66;
  assign T66 = io_req_bits_tag_match ^ 1'h1;
  assign T67 = io_replay_ready & T68;
  assign T68 = state == 4'h8;
  assign T69 = io_meta_read_ready ^ 1'h1;
  assign T70 = T75 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T74 | T73;
  assign T73 = io_req_bits_cmd == 5'h3;
  assign T74 = io_req_bits_cmd == 5'h2;
  assign T75 = T117 | T76;
  assign T76 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T77;
  assign T77 = T110 | T78;
  assign T78 = T107 & T79;
  assign T79 = cmd_requires_second_acquire ^ 1'h1;
  assign cmd_requires_second_acquire = T96 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T87 | T82;
  assign T82 = req_cmd == 5'h6;
  assign T83 = T60 ? io_req_bits_cmd : T84;
  assign T84 = T85 ? io_req_bits_cmd : req_cmd;
  assign T85 = T86 & cmd_requires_second_acquire;
  assign T86 = io_req_sec_val & io_req_sec_rdy;
  assign T87 = T89 | T88;
  assign T88 = req_cmd == 5'h3;
  assign T89 = T93 | T90;
  assign T90 = T92 | T91;
  assign T91 = req_cmd == 5'h4;
  assign T92 = req_cmd[2'h3:2'h3];
  assign T93 = T95 | T94;
  assign T94 = req_cmd == 5'h7;
  assign T95 = req_cmd == 5'h1;
  assign T96 = T98 | T97;
  assign T97 = io_req_bits_cmd == 5'h6;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h3;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3:2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign T107 = T109 | T108;
  assign T108 = 4'h5 == state;
  assign T109 = 4'h4 == state;
  assign T110 = T112 | T111;
  assign T111 = 4'h3 == state;
  assign T112 = T114 | T113;
  assign T113 = 4'h2 == state;
  assign T114 = 4'h1 == state;
  assign idx_match = req_idx == T115;
  assign T115 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T116 = T60 ? io_req_bits_addr : req_addr;
  assign T117 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T118;
  assign T118 = T132 | T119;
  assign T119 = T126 & T120;
  assign T120 = meta_hazard == 2'h0;
  assign T218 = reset ? 2'h0 : T121;
  assign T121 = T125 ? 2'h1 : T122;
  assign T122 = T124 ? T123 : meta_hazard;
  assign T123 = meta_hazard + 2'h1;
  assign T124 = meta_hazard != 2'h0;
  assign T125 = io_meta_write_ready & io_meta_write_valid;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T129 | T128;
  assign T128 = 4'h3 == state;
  assign T129 = T131 | T130;
  assign T130 = 4'h2 == state;
  assign T131 = 4'h1 == state;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T60 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_data = T134;
  assign T134 = 128'h0;
  assign io_wb_req_bits_voluntary = T135;
  assign T135 = 1'h1;
  assign io_wb_req_bits_r_type = T136;
  assign T136 = T137;
  assign T137 = T138 ? 3'h0 : 3'h3;
  assign T138 = 2'h3 == req_old_meta_coh_state;
  assign T139 = T60 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign io_wb_req_bits_client_xact_id = T140;
  assign T140 = 2'h1;
  assign io_wb_req_bits_addr_block = T141;
  assign T141 = T142;
  assign T142 = {req_old_meta_tag, req_idx};
  assign T143 = T60 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_bits_addr_beat = T144;
  assign T144 = 2'h0;
  assign io_wb_req_valid = T145;
  assign T145 = state == 4'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_cmd = T146;
  assign T146 = T69 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T219;
  assign T219 = {8'h0, T147};
  assign T147 = T148;
  assign T148 = {io_tag, T149};
  assign T149 = {req_idx, T150};
  assign T150 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_valid = T151;
  assign T151 = T152 & rpq_io_deq_valid;
  assign T152 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T153;
  assign T153 = T182 ? T181 : new_coh_state_state;
  assign T154 = 2'h0;
  assign T220 = reset ? T154 : T155;
  assign T155 = T38 ? coh_on_hit_state : T156;
  assign T156 = T172 ? coh_on_grant_state : new_coh_state_state;
  assign coh_on_grant_state = T157;
  assign T157 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T158;
  assign T158 = T171 ? 2'h1 : T159;
  assign T159 = T170 ? T162 : T160;
  assign T160 = T161 ? 2'h3 : 2'h0;
  assign T161 = io_mem_grant_bits_g_type == 4'h2;
  assign T162 = T163 ? 2'h3 : 2'h2;
  assign T163 = T167 | T164;
  assign T164 = T166 | T165;
  assign T165 = req_cmd == 5'h4;
  assign T166 = req_cmd[2'h3:2'h3];
  assign T167 = T169 | T168;
  assign T168 = req_cmd == 5'h7;
  assign T169 = req_cmd == 5'h1;
  assign T170 = io_mem_grant_bits_g_type == 4'h1;
  assign T171 = io_mem_grant_bits_g_type == 4'h0;
  assign T172 = T31 & io_mem_grant_valid;
  assign coh_on_hit_state = T173;
  assign T173 = T174 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T174 = T178 | T175;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h4;
  assign T177 = io_req_bits_cmd[2'h3:2'h3];
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h7;
  assign T180 = io_req_bits_cmd == 5'h1;
  assign T181 = 2'h0;
  assign T182 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T183;
  assign T183 = T185 | T184;
  assign T184 = state == 4'h3;
  assign T185 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T186;
  assign T186 = state == 4'h8;
  assign io_refill_addr = T187;
  assign T187 = T188 << 3'h4;
  assign T188 = {req_idx, refill_cnt};
  assign io_refill_way_en = req_way_en;
  assign io_mem_req_bits_data = T189;
  assign T189 = 128'h0;
  assign io_mem_req_bits_union = T190;
  assign T190 = T221;
  assign T221 = {11'h0, T191};
  assign T191 = {req_cmd, 1'h1};
  assign io_mem_req_bits_a_type = T192;
  assign T192 = T222;
  assign T222 = {2'h0, T193};
  assign T193 = T195 | T194;
  assign T194 = req_cmd == 5'h6;
  assign T195 = T197 | T196;
  assign T196 = req_cmd == 5'h3;
  assign T197 = T201 | T198;
  assign T198 = T200 | T199;
  assign T199 = req_cmd == 5'h4;
  assign T200 = req_cmd[2'h3:2'h3];
  assign T201 = T203 | T202;
  assign T202 = req_cmd == 5'h7;
  assign T203 = req_cmd == 5'h1;
  assign io_mem_req_bits_is_builtin_type = T204;
  assign T204 = 1'h0;
  assign io_mem_req_bits_addr_beat = T205;
  assign T205 = 2'h0;
  assign io_mem_req_bits_client_xact_id = T206;
  assign T206 = 2'h1;
  assign io_mem_req_bits_addr_block = T207;
  assign T207 = T208;
  assign T208 = T209;
  assign T209 = {io_tag, req_idx};
  assign io_mem_req_valid = T210;
  assign T210 = state == 4'h4;
  assign io_tag = T223;
  assign T223 = T211[5'h13:1'h0];
  assign T211 = req_addr >> 4'hc;
  assign io_idx_match = T212;
  assign T212 = T213 & idx_match;
  assign T213 = state != 4'h0;
  assign io_req_sec_rdy = T214;
  assign T214 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T215;
  assign T215 = state == 4'h0;
  Queue_14 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T70 ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T65) begin
      state <= T63;
    end else if(T61) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T24;
    end
    if(T60) begin
      req_cmd <= io_req_bits_cmd;
    end else if(T85) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T60) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T125) begin
      meta_hazard <= 2'h1;
    end else if(T124) begin
      meta_hazard <= T123;
    end
    if(T60) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T60) begin
      req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
    end
    if(T60) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(reset) begin
      new_coh_state_state <= T154;
    end else if(T38) begin
      new_coh_state_state <= coh_on_hit_state;
    end else if(T172) begin
      new_coh_state_state <= coh_on_grant_state;
    end
  end
endmodule

module Arbiter_9(
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire chosen;


  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits = io_in_0_bits;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
endmodule

module Arbiter_10(
    output io_in_0_ready,
    input  io_in_0_valid,
    input [39:0] io_in_0_bits_addr,
    input [8:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [2:0] io_in_0_bits_typ,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_nack,
    input  io_in_0_bits_replay,
    input  io_in_0_bits_has_data,
    input [63:0] io_in_0_bits_data_word_bypass,
    input [63:0] io_in_0_bits_store_data,
    input  io_out_ready,
    output io_out_valid,
    output[39:0] io_out_bits_addr,
    output[8:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[2:0] io_out_bits_typ,
    output[63:0] io_out_bits_data,
    output io_out_bits_nack,
    output io_out_bits_replay,
    output io_out_bits_has_data,
    output[63:0] io_out_bits_data_word_bypass,
    output[63:0] io_out_bits_store_data,
    output io_chosen
);

  wire chosen;


  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits_store_data = io_in_0_bits_store_data;
  assign io_out_bits_data_word_bypass = io_in_0_bits_data_word_bypass;
  assign io_out_bits_has_data = io_in_0_bits_has_data;
  assign io_out_bits_replay = io_in_0_bits_replay;
  assign io_out_bits_nack = io_in_0_bits_nack;
  assign io_out_bits_data = io_in_0_bits_data;
  assign io_out_bits_typ = io_in_0_bits_typ;
  assign io_out_bits_cmd = io_in_0_bits_cmd;
  assign io_out_bits_tag = io_in_0_bits_tag;
  assign io_out_bits_addr = io_in_0_bits_addr;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
endmodule

module IOMSHR(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [39:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [63:0] io_req_bits_data,
    input  io_acquire_ready,
    output io_acquire_valid,
    output[25:0] io_acquire_bits_addr_block,
    output[1:0] io_acquire_bits_client_xact_id,
    output[1:0] io_acquire_bits_addr_beat,
    output io_acquire_bits_is_builtin_type,
    output[2:0] io_acquire_bits_a_type,
    output[16:0] io_acquire_bits_union,
    output[127:0] io_acquire_bits_data,
    input  io_grant_valid,
    input [1:0] io_grant_bits_addr_beat,
    input [1:0] io_grant_bits_client_xact_id,
    input [3:0] io_grant_bits_manager_xact_id,
    input  io_grant_bits_is_builtin_type,
    input [3:0] io_grant_bits_g_type,
    input [127:0] io_grant_bits_data,
    input  io_resp_ready,
    output io_resp_valid,
    output[39:0] io_resp_bits_addr,
    output[8:0] io_resp_bits_tag,
    output[4:0] io_resp_bits_cmd,
    output[2:0] io_resp_bits_typ,
    output[63:0] io_resp_bits_data,
    output io_resp_bits_nack,
    output io_resp_bits_replay,
    output io_resp_bits_has_data,
    //output[63:0] io_resp_bits_data_word_bypass
    output[63:0] io_resp_bits_store_data
);

  reg [63:0] req_data;
  wire[63:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg [4:0] req_cmd;
  wire[4:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[63:0] T12;
  wire[63:0] T156;
  wire req_cmd_sc;
  wire[63:0] T13;
  wire[7:0] T14;
  wire[7:0] T15;
  wire[7:0] T16;
  wire[63:0] T17;
  wire[15:0] T18;
  wire[15:0] T19;
  wire[63:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  reg [63:0] grant_word;
  wire[63:0] T23;
  wire[63:0] T24;
  wire[127:0] T25;
  wire[6:0] T26;
  wire T27;
  reg [39:0] req_addr;
  wire[39:0] T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg [1:0] state;
  wire[1:0] T157;
  wire[1:0] T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[31:0] T50;
  wire T51;
  wire[31:0] T52;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T158;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  reg [2:0] req_typ;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[15:0] T68;
  wire T69;
  wire[47:0] T70;
  wire[47:0] T71;
  wire[47:0] T72;
  wire[47:0] T159;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire T79;
  wire[55:0] T80;
  wire[55:0] T81;
  wire[55:0] T82;
  wire[55:0] T160;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  reg [8:0] req_tag;
  wire[8:0] T89;
  wire T90;
  wire[127:0] T91;
  wire[127:0] beat_data;
  wire[63:0] T92;
  wire[63:0] T93;
  wire[63:0] T94;
  wire[63:0] T95;
  wire[31:0] T96;
  wire T97;
  wire T98;
  wire T99;
  wire[63:0] T100;
  wire[31:0] T101;
  wire[15:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire[63:0] T106;
  wire[31:0] T107;
  wire[15:0] T108;
  wire[7:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[16:0] T113;
  wire[16:0] T161;
  wire[26:0] T114;
  wire[25:0] union;
  wire[25:0] beat_mask;
  wire[3:0] T115;
  wire beat_offset;
  wire[10:0] T116;
  wire[10:0] T117;
  wire[10:0] T118;
  wire[10:0] T119;
  wire[2:0] T120;
  wire T121;
  wire[10:0] T162;
  wire[8:0] T122;
  wire[2:0] T123;
  wire[1:0] T124;
  wire[10:0] T163;
  wire[7:0] T125;
  wire[2:0] T126;
  wire[25:0] T164;
  wire[11:0] T127;
  wire[7:0] T128;
  wire[3:0] addr_byte;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire[2:0] T138;
  wire[2:0] a_type;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire[1:0] T149;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[25:0] T152;
  wire[25:0] T153;
  wire T154;
  wire T155;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_data = {2{$random}};
    req_cmd = {1{$random}};
    grant_word = {2{$random}};
    req_addr = {2{$random}};
    state = {1{$random}};
    req_typ = {1{$random}};
    req_tag = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_resp_bits_data_word_bypass = {2{$random}};
// synthesis translate_on
`endif
  assign io_resp_bits_store_data = req_data;
  assign T0 = T1 ? io_req_bits_data : req_data;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_has_data = T2;
  assign T2 = T7 | T3;
  assign T3 = T6 | T4;
  assign T4 = req_cmd == 5'h4;
  assign T5 = T1 ? io_req_bits_cmd : req_cmd;
  assign T6 = req_cmd[2'h3:2'h3];
  assign T7 = T9 | T8;
  assign T8 = req_cmd == 5'h7;
  assign T9 = T11 | T10;
  assign T10 = req_cmd == 5'h6;
  assign T11 = req_cmd == 5'h0;
  assign io_resp_bits_replay = io_resp_valid;
  assign io_resp_bits_nack = 1'h0;
  assign io_resp_bits_data = T12;
  assign T12 = T13 | T156;
  assign T156 = {63'h0, req_cmd_sc};
  assign req_cmd_sc = req_cmd == 5'h7;
  assign T13 = {T80, T14};
  assign T14 = req_cmd_sc ? 8'h0 : T15;
  assign T15 = T79 ? T78 : T16;
  assign T16 = T17[3'h7:1'h0];
  assign T17 = {T70, T18};
  assign T18 = T69 ? T68 : T19;
  assign T19 = T20[4'hf:1'h0];
  assign T20 = {T52, T21};
  assign T21 = T51 ? T50 : T22;
  assign T22 = grant_word[5'h1f:1'h0];
  assign T23 = T29 ? T24 : grant_word;
  assign T24 = T25[6'h3f:1'h0];
  assign T25 = io_grant_bits_data >> T26;
  assign T26 = {T27, 6'h0};
  assign T27 = req_addr[2'h3:2'h3];
  assign T28 = T1 ? io_req_bits_addr : req_addr;
  assign T29 = T39 & T30;
  assign T30 = T34 | T31;
  assign T31 = T33 | T32;
  assign T32 = req_cmd == 5'h4;
  assign T33 = req_cmd[2'h3:2'h3];
  assign T34 = T36 | T35;
  assign T35 = req_cmd == 5'h7;
  assign T36 = T38 | T37;
  assign T37 = req_cmd == 5'h6;
  assign T38 = req_cmd == 5'h0;
  assign T39 = T40 & io_grant_valid;
  assign T40 = state == 2'h2;
  assign T157 = reset ? 2'h0 : T41;
  assign T41 = T49 ? 2'h0 : T42;
  assign T42 = T47 ? 2'h0 : T43;
  assign T43 = T29 ? 2'h3 : T44;
  assign T44 = T46 ? 2'h2 : T45;
  assign T45 = T1 ? 2'h1 : state;
  assign T46 = io_acquire_ready & io_acquire_valid;
  assign T47 = T39 & T48;
  assign T48 = T30 ^ 1'h1;
  assign T49 = io_resp_ready & io_resp_valid;
  assign T50 = grant_word[6'h3f:6'h20];
  assign T51 = req_addr[2'h2:2'h2];
  assign T52 = T65 ? T54 : T53;
  assign T53 = grant_word[6'h3f:6'h20];
  assign T54 = 32'h0 - T158;
  assign T158 = {31'h0, T55};
  assign T55 = T57 & T56;
  assign T56 = T21[5'h1f:5'h1f];
  assign T57 = T60 | T58;
  assign T58 = req_typ == 3'h3;
  assign T59 = T1 ? io_req_bits_typ : req_typ;
  assign T60 = T62 | T61;
  assign T61 = req_typ == 3'h2;
  assign T62 = T64 | T63;
  assign T63 = req_typ == 3'h1;
  assign T64 = req_typ == 3'h0;
  assign T65 = T67 | T66;
  assign T66 = req_typ == 3'h6;
  assign T67 = req_typ == 3'h2;
  assign T68 = T20[5'h1f:5'h10];
  assign T69 = req_addr[1'h1:1'h1];
  assign T70 = T75 ? T72 : T71;
  assign T71 = T20[6'h3f:5'h10];
  assign T72 = 48'h0 - T159;
  assign T159 = {47'h0, T73};
  assign T73 = T57 & T74;
  assign T74 = T18[4'hf:4'hf];
  assign T75 = T77 | T76;
  assign T76 = req_typ == 3'h5;
  assign T77 = req_typ == 3'h1;
  assign T78 = T17[4'hf:4'h8];
  assign T79 = req_addr[1'h0:1'h0];
  assign T80 = T85 ? T82 : T81;
  assign T81 = T17[6'h3f:4'h8];
  assign T82 = 56'h0 - T160;
  assign T160 = {55'h0, T83};
  assign T83 = T57 & T84;
  assign T84 = T14[3'h7:3'h7];
  assign T85 = req_cmd_sc | T86;
  assign T86 = T88 | T87;
  assign T87 = req_typ == 3'h4;
  assign T88 = req_typ == 3'h0;
  assign io_resp_bits_typ = req_typ;
  assign io_resp_bits_cmd = req_cmd;
  assign io_resp_bits_tag = req_tag;
  assign T89 = T1 ? io_req_bits_tag : req_tag;
  assign io_resp_bits_addr = req_addr;
  assign io_resp_valid = T90;
  assign T90 = state == 2'h3;
  assign io_acquire_bits_data = T91;
  assign T91 = beat_data;
  assign beat_data = {T92, T92};
  assign T92 = T110 ? T106 : T93;
  assign T93 = T103 ? T100 : T94;
  assign T94 = T97 ? T95 : req_data;
  assign T95 = {T96, T96};
  assign T96 = req_data[5'h1f:1'h0];
  assign T97 = T99 | T98;
  assign T98 = req_typ == 3'h6;
  assign T99 = req_typ == 3'h2;
  assign T100 = {T101, T101};
  assign T101 = {T102, T102};
  assign T102 = req_data[4'hf:1'h0];
  assign T103 = T105 | T104;
  assign T104 = req_typ == 3'h5;
  assign T105 = req_typ == 3'h1;
  assign T106 = {T107, T107};
  assign T107 = {T108, T108};
  assign T108 = {T109, T109};
  assign T109 = req_data[3'h7:1'h0];
  assign T110 = T112 | T111;
  assign T111 = req_typ == 3'h4;
  assign T112 = req_typ == 3'h0;
  assign io_acquire_bits_union = T113;
  assign T113 = T161;
  assign T161 = T114[5'h10:1'h0];
  assign T114 = {union, 1'h0};
  assign union = T129 ? T164 : beat_mask;
  assign beat_mask = T116 << T115;
  assign T115 = {beat_offset, 3'h0};
  assign beat_offset = req_addr[2'h3:2'h3];
  assign T116 = T110 ? T163 : T117;
  assign T117 = T103 ? T162 : T118;
  assign T118 = T97 ? T119 : 11'hff;
  assign T119 = 4'hf << T120;
  assign T120 = {T121, 2'h0};
  assign T121 = req_addr[2'h2:2'h2];
  assign T162 = {2'h0, T122};
  assign T122 = 2'h3 << T123;
  assign T123 = {T124, 1'h0};
  assign T124 = req_addr[2'h2:1'h1];
  assign T163 = {3'h0, T125};
  assign T125 = 1'h1 << T126;
  assign T126 = req_addr[2'h2:1'h0];
  assign T164 = {14'h0, T127};
  assign T127 = {addr_byte, T128};
  assign T128 = {req_typ, 5'h0};
  assign addr_byte = req_addr[2'h3:1'h0];
  assign T129 = T133 | T130;
  assign T130 = T132 | T131;
  assign T131 = req_cmd == 5'h4;
  assign T132 = req_cmd[2'h3:2'h3];
  assign T133 = T135 | T134;
  assign T134 = req_cmd == 5'h7;
  assign T135 = T137 | T136;
  assign T136 = req_cmd == 5'h6;
  assign T137 = req_cmd == 5'h0;
  assign io_acquire_bits_a_type = T138;
  assign T138 = a_type;
  assign a_type = T139 ? 3'h0 : 3'h2;
  assign T139 = T143 | T140;
  assign T140 = T142 | T141;
  assign T141 = req_cmd == 5'h4;
  assign T142 = req_cmd[2'h3:2'h3];
  assign T143 = T145 | T144;
  assign T144 = req_cmd == 5'h7;
  assign T145 = T147 | T146;
  assign T146 = req_cmd == 5'h6;
  assign T147 = req_cmd == 5'h0;
  assign io_acquire_bits_is_builtin_type = T148;
  assign T148 = 1'h1;
  assign io_acquire_bits_addr_beat = T149;
  assign T149 = T150;
  assign T150 = req_addr[3'h5:3'h4];
  assign io_acquire_bits_client_xact_id = T151;
  assign T151 = 2'h2;
  assign io_acquire_bits_addr_block = T152;
  assign T152 = T153;
  assign T153 = req_addr[5'h1f:3'h6];
  assign io_acquire_valid = T154;
  assign T154 = state == 2'h1;
  assign io_req_ready = T155;
  assign T155 = state == 2'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_data <= io_req_bits_data;
    end
    if(T1) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T29) begin
      grant_word <= T24;
    end
    if(T1) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T49) begin
      state <= 2'h0;
    end else if(T47) begin
      state <= 2'h0;
    end else if(T29) begin
      state <= 2'h3;
    end else if(T46) begin
      state <= 2'h2;
    end else if(T1) begin
      state <= 2'h1;
    end
    if(T1) begin
      req_typ <= io_req_bits_typ;
    end
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [39:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [63:0] io_req_bits_data,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    input  io_resp_ready,
    output io_resp_valid,
    output[39:0] io_resp_bits_addr,
    output[8:0] io_resp_bits_tag,
    output[4:0] io_resp_bits_cmd,
    output[2:0] io_resp_bits_typ,
    output[63:0] io_resp_bits_data,
    output io_resp_bits_nack,
    output io_resp_bits_replay,
    output io_resp_bits_has_data,
    output[63:0] io_resp_bits_data_word_bypass,
    output[63:0] io_resp_bits_store_data,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output[127:0] io_mem_req_bits_data,
    output[3:0] io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[8:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[63:0] io_replay_bits_data,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_wb_req_bits_voluntary,
    output[127:0] io_wb_req_bits_data,
    output[3:0] io_wb_req_bits_way_en,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[4:0] T86;
  wire[4:0] T87;
  wire[4:0] T88;
  wire[4:0] T89;
  wire[4:0] T90;
  wire[4:0] T91;
  wire[4:0] T92;
  wire[4:0] T93;
  wire[4:0] T94;
  wire[4:0] T95;
  wire[4:0] T96;
  wire[4:0] T97;
  wire[4:0] T98;
  wire[4:0] T99;
  wire[4:0] T100;
  wire[4:0] T101;
  wire T102;
  wire[16:0] T4;
  wire[16:0] T5;
  reg [16:0] sdq_val;
  wire[16:0] T103;
  wire[31:0] T104;
  wire[31:0] T6;
  wire[31:0] T105;
  wire[31:0] T7;
  wire[31:0] T106;
  wire[16:0] T8;
  wire[16:0] T9;
  wire[16:0] T10;
  wire[16:0] T11;
  wire[16:0] T12;
  wire[16:0] T13;
  wire[16:0] T14;
  wire[16:0] T15;
  wire[16:0] T16;
  wire[16:0] T17;
  wire[16:0] T18;
  wire[16:0] T19;
  wire[16:0] T20;
  wire[16:0] T21;
  wire[16:0] T22;
  wire[16:0] T23;
  wire[16:0] T24;
  wire[16:0] T25;
  wire T26;
  wire[16:0] T27;
  wire[16:0] T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[31:0] T45;
  wire[31:0] T46;
  wire[31:0] T47;
  wire[31:0] T107;
  wire[16:0] T48;
  wire[16:0] T108;
  wire free_sdq;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[31:0] T57;
  wire[31:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T58;
  wire tag_match;
  wire[27:0] T59;
  wire[27:0] T125;
  wire[19:0] T60;
  wire[19:0] T61;
  wire[19:0] tagList_1;
  wire idxMatch_1;
  wire[19:0] T62;
  wire[19:0] tagList_0;
  wire idxMatch_0;
  wire T63;
  wire sdq_rdy;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire[63:0] T79;
  reg [63:0] sdq [16:0];
  wire[63:0] T80;
  reg [4:0] R81;
  wire[4:0] T82;
  wire[11:0] T83;
  wire[11:0] refillMux_0_addr;
  wire[11:0] refillMux_1_addr;
  wire T84;
  wire T126;
  wire[3:0] T85;
  wire[3:0] refillMux_0_way_en;
  wire[3:0] refillMux_1_way_en;
  wire idx_match;
  wire meta_read_arb_io_in_1_ready;
  wire meta_read_arb_io_in_0_ready;
  wire meta_read_arb_io_out_valid;
  wire[5:0] meta_read_arb_io_out_bits_idx;
  wire[19:0] meta_read_arb_io_out_bits_tag;
  wire meta_write_arb_io_in_1_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_write_arb_io_out_valid;
  wire[5:0] meta_write_arb_io_out_bits_idx;
  wire[3:0] meta_write_arb_io_out_bits_way_en;
  wire[19:0] meta_write_arb_io_out_bits_data_tag;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire mem_req_arb_io_in_2_ready;
  wire mem_req_arb_io_in_1_ready;
  wire mem_req_arb_io_in_0_ready;
  wire mem_req_arb_io_out_valid;
  wire[25:0] mem_req_arb_io_out_bits_addr_block;
  wire[1:0] mem_req_arb_io_out_bits_client_xact_id;
  wire[1:0] mem_req_arb_io_out_bits_addr_beat;
  wire mem_req_arb_io_out_bits_is_builtin_type;
  wire[2:0] mem_req_arb_io_out_bits_a_type;
  wire[16:0] mem_req_arb_io_out_bits_union;
  wire[127:0] mem_req_arb_io_out_bits_data;
  wire wb_req_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire wb_req_arb_io_out_valid;
  wire[1:0] wb_req_arb_io_out_bits_addr_beat;
  wire[25:0] wb_req_arb_io_out_bits_addr_block;
  wire[1:0] wb_req_arb_io_out_bits_client_xact_id;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire wb_req_arb_io_out_bits_voluntary;
  wire[127:0] wb_req_arb_io_out_bits_data;
  wire[3:0] wb_req_arb_io_out_bits_way_en;
  wire replay_arb_io_in_1_ready;
  wire replay_arb_io_in_0_ready;
  wire replay_arb_io_out_valid;
  wire[39:0] replay_arb_io_out_bits_addr;
  wire[8:0] replay_arb_io_out_bits_tag;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[2:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_kill;
  wire replay_arb_io_out_bits_phys;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire mmio_alloc_arb_io_in_0_ready;
  wire resp_arb_io_in_0_ready;
  wire resp_arb_io_out_valid;
  wire[39:0] resp_arb_io_out_bits_addr;
  wire[8:0] resp_arb_io_out_bits_tag;
  wire[4:0] resp_arb_io_out_bits_cmd;
  wire[2:0] resp_arb_io_out_bits_typ;
  wire[63:0] resp_arb_io_out_bits_data;
  wire resp_arb_io_out_bits_nack;
  wire resp_arb_io_out_bits_replay;
  wire resp_arb_io_out_bits_has_data;
  wire[63:0] resp_arb_io_out_bits_data_word_bypass;
  wire[63:0] resp_arb_io_out_bits_store_data;
  wire IOMSHR_io_req_ready;
  wire IOMSHR_io_acquire_valid;
  wire[25:0] IOMSHR_io_acquire_bits_addr_block;
  wire[1:0] IOMSHR_io_acquire_bits_client_xact_id;
  wire[1:0] IOMSHR_io_acquire_bits_addr_beat;
  wire IOMSHR_io_acquire_bits_is_builtin_type;
  wire[2:0] IOMSHR_io_acquire_bits_a_type;
  wire[16:0] IOMSHR_io_acquire_bits_union;
  wire[127:0] IOMSHR_io_acquire_bits_data;
  wire IOMSHR_io_resp_valid;
  wire[39:0] IOMSHR_io_resp_bits_addr;
  wire[8:0] IOMSHR_io_resp_bits_tag;
  wire[4:0] IOMSHR_io_resp_bits_cmd;
  wire[2:0] IOMSHR_io_resp_bits_typ;
  wire[63:0] IOMSHR_io_resp_bits_data;
  wire IOMSHR_io_resp_bits_nack;
  wire IOMSHR_io_resp_bits_replay;
  wire IOMSHR_io_resp_bits_has_data;
  wire[63:0] IOMSHR_io_resp_bits_store_data;
  wire MSHR_io_req_pri_rdy;
  wire MSHR_io_idx_match;
  wire[19:0] MSHR_io_tag;
  wire MSHR_io_mem_req_valid;
  wire[25:0] MSHR_io_mem_req_bits_addr_block;
  wire[1:0] MSHR_io_mem_req_bits_client_xact_id;
  wire[1:0] MSHR_io_mem_req_bits_addr_beat;
  wire MSHR_io_mem_req_bits_is_builtin_type;
  wire[2:0] MSHR_io_mem_req_bits_a_type;
  wire[16:0] MSHR_io_mem_req_bits_union;
  wire[127:0] MSHR_io_mem_req_bits_data;
  wire[3:0] MSHR_io_refill_way_en;
  wire[11:0] MSHR_io_refill_addr;
  wire MSHR_io_meta_read_valid;
  wire[5:0] MSHR_io_meta_read_bits_idx;
  wire[19:0] MSHR_io_meta_read_bits_tag;
  wire MSHR_io_meta_write_valid;
  wire[5:0] MSHR_io_meta_write_bits_idx;
  wire[3:0] MSHR_io_meta_write_bits_way_en;
  wire[19:0] MSHR_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_io_meta_write_bits_data_coh_state;
  wire MSHR_io_replay_valid;
  wire[39:0] MSHR_io_replay_bits_addr;
  wire[8:0] MSHR_io_replay_bits_tag;
  wire[4:0] MSHR_io_replay_bits_cmd;
  wire[2:0] MSHR_io_replay_bits_typ;
  wire MSHR_io_replay_bits_kill;
  wire MSHR_io_replay_bits_phys;
  wire[4:0] MSHR_io_replay_bits_sdq_id;
  wire MSHR_io_wb_req_valid;
  wire[1:0] MSHR_io_wb_req_bits_addr_beat;
  wire[25:0] MSHR_io_wb_req_bits_addr_block;
  wire[1:0] MSHR_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_io_wb_req_bits_r_type;
  wire MSHR_io_wb_req_bits_voluntary;
  wire[127:0] MSHR_io_wb_req_bits_data;
  wire[3:0] MSHR_io_wb_req_bits_way_en;
  wire MSHR_io_probe_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire MSHR_1_io_idx_match;
  wire[19:0] MSHR_1_io_tag;
  wire MSHR_1_io_mem_req_valid;
  wire[25:0] MSHR_1_io_mem_req_bits_addr_block;
  wire[1:0] MSHR_1_io_mem_req_bits_client_xact_id;
  wire[1:0] MSHR_1_io_mem_req_bits_addr_beat;
  wire MSHR_1_io_mem_req_bits_is_builtin_type;
  wire[2:0] MSHR_1_io_mem_req_bits_a_type;
  wire[16:0] MSHR_1_io_mem_req_bits_union;
  wire[127:0] MSHR_1_io_mem_req_bits_data;
  wire[3:0] MSHR_1_io_refill_way_en;
  wire[11:0] MSHR_1_io_refill_addr;
  wire MSHR_1_io_meta_read_valid;
  wire[5:0] MSHR_1_io_meta_read_bits_idx;
  wire[19:0] MSHR_1_io_meta_read_bits_tag;
  wire MSHR_1_io_meta_write_valid;
  wire[5:0] MSHR_1_io_meta_write_bits_idx;
  wire[3:0] MSHR_1_io_meta_write_bits_way_en;
  wire[19:0] MSHR_1_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire MSHR_1_io_replay_valid;
  wire[39:0] MSHR_1_io_replay_bits_addr;
  wire[8:0] MSHR_1_io_replay_bits_tag;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[2:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_kill;
  wire MSHR_1_io_replay_bits_phys;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire MSHR_1_io_wb_req_valid;
  wire[1:0] MSHR_1_io_wb_req_bits_addr_beat;
  wire[25:0] MSHR_1_io_wb_req_bits_addr_block;
  wire[1:0] MSHR_1_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire MSHR_1_io_wb_req_bits_voluntary;
  wire[127:0] MSHR_1_io_wb_req_bits_data;
  wire[3:0] MSHR_1_io_wb_req_bits_way_en;
  wire MSHR_1_io_probe_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R81 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_mem_grant_valid & T1;
  assign T1 = io_mem_grant_bits_client_xact_id == 2'h2;
  assign T2 = io_mem_grant_valid & T3;
  assign T3 = io_mem_grant_bits_client_xact_id == 2'h1;
  assign T86 = T124 ? 1'h0 : T87;
  assign T87 = T123 ? 1'h1 : T88;
  assign T88 = T122 ? 2'h2 : T89;
  assign T89 = T121 ? 2'h3 : T90;
  assign T90 = T120 ? 3'h4 : T91;
  assign T91 = T119 ? 3'h5 : T92;
  assign T92 = T118 ? 3'h6 : T93;
  assign T93 = T117 ? 3'h7 : T94;
  assign T94 = T116 ? 4'h8 : T95;
  assign T95 = T115 ? 4'h9 : T96;
  assign T96 = T114 ? 4'ha : T97;
  assign T97 = T113 ? 4'hb : T98;
  assign T98 = T112 ? 4'hc : T99;
  assign T99 = T111 ? 4'hd : T100;
  assign T100 = T110 ? 4'he : T101;
  assign T101 = T102 ? 4'hf : 5'h10;
  assign T102 = T4[4'hf:4'hf];
  assign T4 = ~ T5;
  assign T5 = sdq_val[5'h10:1'h0];
  assign T103 = T104[5'h10:1'h0];
  assign T104 = reset ? 32'h0 : T6;
  assign T6 = io_replay_valid ? T7 : T105;
  assign T105 = {15'h0, sdq_val};
  assign T7 = T45 | T106;
  assign T106 = {15'h0, T8};
  assign T8 = T9 & 17'h0;
  assign T9 = T44 ? 17'h1 : T10;
  assign T10 = T43 ? 17'h2 : T11;
  assign T11 = T42 ? 17'h4 : T12;
  assign T12 = T41 ? 17'h8 : T13;
  assign T13 = T40 ? 17'h10 : T14;
  assign T14 = T39 ? 17'h20 : T15;
  assign T15 = T38 ? 17'h40 : T16;
  assign T16 = T37 ? 17'h80 : T17;
  assign T17 = T36 ? 17'h100 : T18;
  assign T18 = T35 ? 17'h200 : T19;
  assign T19 = T34 ? 17'h400 : T20;
  assign T20 = T33 ? 17'h800 : T21;
  assign T21 = T32 ? 17'h1000 : T22;
  assign T22 = T31 ? 17'h2000 : T23;
  assign T23 = T30 ? 17'h4000 : T24;
  assign T24 = T29 ? 17'h8000 : T25;
  assign T25 = T26 ? 17'h10000 : 17'h0;
  assign T26 = T27[5'h10:5'h10];
  assign T27 = ~ T28;
  assign T28 = sdq_val[5'h10:1'h0];
  assign T29 = T27[4'hf:4'hf];
  assign T30 = T27[4'he:4'he];
  assign T31 = T27[4'hd:4'hd];
  assign T32 = T27[4'hc:4'hc];
  assign T33 = T27[4'hb:4'hb];
  assign T34 = T27[4'ha:4'ha];
  assign T35 = T27[4'h9:4'h9];
  assign T36 = T27[4'h8:4'h8];
  assign T37 = T27[3'h7:3'h7];
  assign T38 = T27[3'h6:3'h6];
  assign T39 = T27[3'h5:3'h5];
  assign T40 = T27[3'h4:3'h4];
  assign T41 = T27[2'h3:2'h3];
  assign T42 = T27[2'h2:2'h2];
  assign T43 = T27[1'h1:1'h1];
  assign T44 = T27[1'h0:1'h0];
  assign T45 = T109 & T46;
  assign T46 = ~ T47;
  assign T47 = T57 & T107;
  assign T107 = {15'h0, T48};
  assign T48 = 17'h0 - T108;
  assign T108 = {16'h0, free_sdq};
  assign free_sdq = T56 & T49;
  assign T49 = T53 | T50;
  assign T50 = T52 | T51;
  assign T51 = io_replay_bits_cmd == 5'h4;
  assign T52 = io_replay_bits_cmd[2'h3:2'h3];
  assign T53 = T55 | T54;
  assign T54 = io_replay_bits_cmd == 5'h7;
  assign T55 = io_replay_bits_cmd == 5'h1;
  assign T56 = io_replay_ready & io_replay_valid;
  assign T57 = 1'h1 << replay_arb_io_out_bits_sdq_id;
  assign T109 = {15'h0, sdq_val};
  assign T110 = T4[4'he:4'he];
  assign T111 = T4[4'hd:4'hd];
  assign T112 = T4[4'hc:4'hc];
  assign T113 = T4[4'hb:4'hb];
  assign T114 = T4[4'ha:4'ha];
  assign T115 = T4[4'h9:4'h9];
  assign T116 = T4[4'h8:4'h8];
  assign T117 = T4[3'h7:3'h7];
  assign T118 = T4[3'h6:3'h6];
  assign T119 = T4[3'h5:3'h5];
  assign T120 = T4[3'h4:3'h4];
  assign T121 = T4[2'h3:2'h3];
  assign T122 = T4[2'h2:2'h2];
  assign T123 = T4[1'h1:1'h1];
  assign T124 = T4[1'h0:1'h0];
  assign T58 = T63 & tag_match;
  assign tag_match = T125 == T59;
  assign T59 = io_req_bits_addr >> 4'hc;
  assign T125 = {8'h0, T60};
  assign T60 = T62 | T61;
  assign T61 = idxMatch_1 ? tagList_1 : 20'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T62 = idxMatch_0 ? tagList_0 : 20'h0;
  assign tagList_0 = MSHR_io_tag;
  assign idxMatch_0 = MSHR_io_idx_match;
  assign T63 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T64 ^ 1'h1;
  assign T64 = sdq_val == 17'h1ffff;
  assign T65 = io_mem_grant_valid & T66;
  assign T66 = io_mem_grant_bits_client_xact_id == 2'h0;
  assign T67 = T68 & tag_match;
  assign T68 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T69;
  assign T69 = T74 ? 1'h0 : T70;
  assign T70 = T73 ? 1'h0 : T71;
  assign T71 = T72 == 1'h0;
  assign T72 = MSHR_io_req_pri_rdy ^ 1'h1;
  assign T73 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign T74 = IOMSHR_io_req_ready ^ 1'h1;
  assign io_probe_rdy = T75;
  assign T75 = T78 ? 1'h0 : T76;
  assign T76 = T77 == 1'h0;
  assign T77 = MSHR_io_probe_rdy ^ 1'h1;
  assign T78 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_data = wb_req_arb_io_out_bits_data;
  assign io_wb_req_bits_voluntary = wb_req_arb_io_out_bits_voluntary;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_addr_block = wb_req_arb_io_out_bits_addr_block;
  assign io_wb_req_bits_addr_beat = wb_req_arb_io_out_bits_addr_beat;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_replay_bits_data = T79;
  assign T79 = sdq[R81];
  assign T82 = free_sdq ? replay_arb_io_out_bits_sdq_id : R81;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_refill_addr = T83;
  assign T83 = T84 ? refillMux_1_addr : refillMux_0_addr;
  assign refillMux_0_addr = MSHR_io_refill_addr;
  assign refillMux_1_addr = MSHR_1_io_refill_addr;
  assign T84 = T126;
  assign T126 = io_mem_grant_bits_client_xact_id[1'h0:1'h0];
  assign io_refill_way_en = T85;
  assign T85 = T84 ? refillMux_1_way_en : refillMux_0_way_en;
  assign refillMux_0_way_en = MSHR_io_refill_way_en;
  assign refillMux_1_way_en = MSHR_1_io_refill_way_en;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_union = mem_req_arb_io_out_bits_union;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_is_builtin_type = mem_req_arb_io_out_bits_is_builtin_type;
  assign io_mem_req_bits_addr_beat = mem_req_arb_io_out_bits_addr_beat;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr_block = mem_req_arb_io_out_bits_addr_block;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign idx_match = MSHR_io_idx_match | MSHR_1_io_idx_match;
  assign io_resp_bits_store_data = resp_arb_io_out_bits_store_data;
  assign io_resp_bits_data_word_bypass = resp_arb_io_out_bits_data_word_bypass;
  assign io_resp_bits_has_data = resp_arb_io_out_bits_has_data;
  assign io_resp_bits_replay = resp_arb_io_out_bits_replay;
  assign io_resp_bits_nack = resp_arb_io_out_bits_nack;
  assign io_resp_bits_data = resp_arb_io_out_bits_data;
  assign io_resp_bits_typ = resp_arb_io_out_bits_typ;
  assign io_resp_bits_cmd = resp_arb_io_out_bits_cmd;
  assign io_resp_bits_tag = resp_arb_io_out_bits_tag;
  assign io_resp_bits_addr = resp_arb_io_out_bits_addr;
  assign io_resp_valid = resp_arb_io_out_valid;
  assign io_req_ready = IOMSHR_io_req_ready;
  Arbiter_6 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_io_meta_read_bits_idx ),
       .io_in_0_bits_tag( MSHR_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  LockingArbiter_1 mem_req_arb(.clk(clk), .reset(reset),
       .io_in_2_ready( mem_req_arb_io_in_2_ready ),
       .io_in_2_valid( IOMSHR_io_acquire_valid ),
       .io_in_2_bits_addr_block( IOMSHR_io_acquire_bits_addr_block ),
       .io_in_2_bits_client_xact_id( IOMSHR_io_acquire_bits_client_xact_id ),
       .io_in_2_bits_addr_beat( IOMSHR_io_acquire_bits_addr_beat ),
       .io_in_2_bits_is_builtin_type( IOMSHR_io_acquire_bits_is_builtin_type ),
       .io_in_2_bits_a_type( IOMSHR_io_acquire_bits_a_type ),
       .io_in_2_bits_union( IOMSHR_io_acquire_bits_union ),
       .io_in_2_bits_data( IOMSHR_io_acquire_bits_data ),
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr_block( MSHR_1_io_mem_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_in_1_bits_addr_beat( MSHR_1_io_mem_req_bits_addr_beat ),
       .io_in_1_bits_is_builtin_type( MSHR_1_io_mem_req_bits_is_builtin_type ),
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_in_1_bits_union( MSHR_1_io_mem_req_bits_union ),
       .io_in_1_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_mem_req_valid ),
       .io_in_0_bits_addr_block( MSHR_io_mem_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( MSHR_io_mem_req_bits_client_xact_id ),
       .io_in_0_bits_addr_beat( MSHR_io_mem_req_bits_addr_beat ),
       .io_in_0_bits_is_builtin_type( MSHR_io_mem_req_bits_is_builtin_type ),
       .io_in_0_bits_a_type( MSHR_io_mem_req_bits_a_type ),
       .io_in_0_bits_union( MSHR_io_mem_req_bits_union ),
       .io_in_0_bits_data( MSHR_io_mem_req_bits_data ),
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr_block( mem_req_arb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( mem_req_arb_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( mem_req_arb_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_union( mem_req_arb_io_out_bits_union ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data )
       //.io_chosen(  )
  );
  Arbiter_4 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_addr_beat( MSHR_1_io_wb_req_bits_addr_beat ),
       .io_in_1_bits_addr_block( MSHR_1_io_wb_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_1_bits_voluntary( MSHR_1_io_wb_req_bits_voluntary ),
       .io_in_1_bits_data( MSHR_1_io_wb_req_bits_data ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_wb_req_valid ),
       .io_in_0_bits_addr_beat( MSHR_io_wb_req_bits_addr_beat ),
       .io_in_0_bits_addr_block( MSHR_io_wb_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( MSHR_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_r_type( MSHR_io_wb_req_bits_r_type ),
       .io_in_0_bits_voluntary( MSHR_io_wb_req_bits_voluntary ),
       .io_in_0_bits_data( MSHR_io_wb_req_bits_data ),
       .io_in_0_bits_way_en( MSHR_io_wb_req_bits_way_en ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_addr_beat( wb_req_arb_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( wb_req_arb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type ),
       .io_out_bits_voluntary( wb_req_arb_io_out_bits_voluntary ),
       .io_out_bits_data( wb_req_arb_io_out_bits_data ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en )
       //.io_chosen(  )
  );
  Arbiter_7 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_replay_valid ),
       .io_in_0_bits_addr( MSHR_io_replay_bits_addr ),
       .io_in_0_bits_tag( MSHR_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_io_replay_bits_cmd ),
       .io_in_0_bits_typ( MSHR_io_replay_bits_typ ),
       .io_in_0_bits_kill( MSHR_io_replay_bits_kill ),
       .io_in_0_bits_phys( MSHR_io_replay_bits_phys ),
       .io_in_0_bits_sdq_id( MSHR_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_8 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( 1'h0 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  MSHR_0 MSHR(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_io_req_pri_rdy ),
       .io_req_sec_val( T67 ),
       //.io_req_sec_rdy(  )
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_sdq_id( T86 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_io_idx_match ),
       .io_tag( MSHR_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( MSHR_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( MSHR_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( MSHR_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_is_builtin_type( MSHR_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( MSHR_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( MSHR_io_mem_req_bits_union ),
       .io_mem_req_bits_data( MSHR_io_mem_req_bits_data ),
       .io_refill_way_en( MSHR_io_refill_way_en ),
       .io_refill_addr( MSHR_io_refill_addr ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_io_replay_valid ),
       .io_replay_bits_addr( MSHR_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_io_replay_bits_cmd ),
       .io_replay_bits_typ( MSHR_io_replay_bits_typ ),
       .io_replay_bits_kill( MSHR_io_replay_bits_kill ),
       .io_replay_bits_phys( MSHR_io_replay_bits_phys ),
       .io_replay_bits_sdq_id( MSHR_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( T65 ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( MSHR_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( MSHR_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( MSHR_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( MSHR_io_wb_req_bits_r_type ),
       .io_wb_req_bits_voluntary( MSHR_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_data( MSHR_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( MSHR_io_wb_req_bits_way_en ),
       .io_probe_rdy( MSHR_io_probe_rdy )
  );
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T58 ),
       //.io_req_sec_rdy(  )
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_sdq_id( T86 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( MSHR_1_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( MSHR_1_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_is_builtin_type( MSHR_1_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( MSHR_1_io_mem_req_bits_union ),
       .io_mem_req_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_refill_way_en( MSHR_1_io_refill_way_en ),
       .io_refill_addr( MSHR_1_io_refill_addr ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( T2 ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( MSHR_1_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( MSHR_1_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_wb_req_bits_voluntary( MSHR_1_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_data( MSHR_1_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );
  Arbiter_9 mmio_alloc_arb(
       .io_in_0_ready( mmio_alloc_arb_io_in_0_ready ),
       .io_in_0_valid( IOMSHR_io_req_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( io_req_valid )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign mmio_alloc_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  Arbiter_10 resp_arb(
       .io_in_0_ready( resp_arb_io_in_0_ready ),
       .io_in_0_valid( IOMSHR_io_resp_valid ),
       .io_in_0_bits_addr( IOMSHR_io_resp_bits_addr ),
       .io_in_0_bits_tag( IOMSHR_io_resp_bits_tag ),
       .io_in_0_bits_cmd( IOMSHR_io_resp_bits_cmd ),
       .io_in_0_bits_typ( IOMSHR_io_resp_bits_typ ),
       .io_in_0_bits_data( IOMSHR_io_resp_bits_data ),
       .io_in_0_bits_nack( IOMSHR_io_resp_bits_nack ),
       .io_in_0_bits_replay( IOMSHR_io_resp_bits_replay ),
       .io_in_0_bits_has_data( IOMSHR_io_resp_bits_has_data ),
       //.io_in_0_bits_data_word_bypass(  )
       .io_in_0_bits_store_data( IOMSHR_io_resp_bits_store_data ),
       .io_out_ready( io_resp_ready ),
       .io_out_valid( resp_arb_io_out_valid ),
       .io_out_bits_addr( resp_arb_io_out_bits_addr ),
       .io_out_bits_tag( resp_arb_io_out_bits_tag ),
       .io_out_bits_cmd( resp_arb_io_out_bits_cmd ),
       .io_out_bits_typ( resp_arb_io_out_bits_typ ),
       .io_out_bits_data( resp_arb_io_out_bits_data ),
       .io_out_bits_nack( resp_arb_io_out_bits_nack ),
       .io_out_bits_replay( resp_arb_io_out_bits_replay ),
       .io_out_bits_has_data( resp_arb_io_out_bits_has_data ),
       .io_out_bits_data_word_bypass( resp_arb_io_out_bits_data_word_bypass ),
       .io_out_bits_store_data( resp_arb_io_out_bits_store_data )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign resp_arb.io_in_0_bits_data_word_bypass = {2{$random}};
// synthesis translate_on
`endif
  IOMSHR IOMSHR(.clk(clk), .reset(reset),
       .io_req_ready( IOMSHR_io_req_ready ),
       .io_req_valid( mmio_alloc_arb_io_in_0_ready ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_data( io_req_bits_data ),
       .io_acquire_ready( mem_req_arb_io_in_2_ready ),
       .io_acquire_valid( IOMSHR_io_acquire_valid ),
       .io_acquire_bits_addr_block( IOMSHR_io_acquire_bits_addr_block ),
       .io_acquire_bits_client_xact_id( IOMSHR_io_acquire_bits_client_xact_id ),
       .io_acquire_bits_addr_beat( IOMSHR_io_acquire_bits_addr_beat ),
       .io_acquire_bits_is_builtin_type( IOMSHR_io_acquire_bits_is_builtin_type ),
       .io_acquire_bits_a_type( IOMSHR_io_acquire_bits_a_type ),
       .io_acquire_bits_union( IOMSHR_io_acquire_bits_union ),
       .io_acquire_bits_data( IOMSHR_io_acquire_bits_data ),
       .io_grant_valid( T0 ),
       .io_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_grant_bits_data( io_mem_grant_bits_data ),
       .io_resp_ready( resp_arb_io_in_0_ready ),
       .io_resp_valid( IOMSHR_io_resp_valid ),
       .io_resp_bits_addr( IOMSHR_io_resp_bits_addr ),
       .io_resp_bits_tag( IOMSHR_io_resp_bits_tag ),
       .io_resp_bits_cmd( IOMSHR_io_resp_bits_cmd ),
       .io_resp_bits_typ( IOMSHR_io_resp_bits_typ ),
       .io_resp_bits_data( IOMSHR_io_resp_bits_data ),
       .io_resp_bits_nack( IOMSHR_io_resp_bits_nack ),
       .io_resp_bits_replay( IOMSHR_io_resp_bits_replay ),
       .io_resp_bits_has_data( IOMSHR_io_resp_bits_has_data ),
       //.io_resp_bits_data_word_bypass(  )
       .io_resp_bits_store_data( IOMSHR_io_resp_bits_store_data )
  );

  always @(posedge clk) begin
    sdq_val <= T103;
    if (1'h0)
      sdq[T86] <= io_req_bits_data;
    if(free_sdq) begin
      R81 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [5:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [5:0] io_write_bits_idx,
    input [3:0] io_write_bits_way_en,
    input [19:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[19:0] io_resp_3_tag,
    output[1:0] io_resp_3_coh_state,
    output[19:0] io_resp_2_tag,
    output[1:0] io_resp_2_coh_state,
    output[19:0] io_resp_1_tag,
    output[1:0] io_resp_1_coh_state,
    output[19:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state
);

  wire[1:0] T0;
  wire[87:0] tags;
  wire[87:0] T1;
  wire[43:0] T2;
  wire[21:0] T3;
  wire[87:0] T4;
  wire[87:0] T5;
  wire[87:0] T6;
  wire[87:0] T7;
  wire[43:0] T8;
  wire[21:0] T9;
  wire[21:0] T48;
  wire T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire rst;
  reg [6:0] rst_cnt;
  wire[6:0] T49;
  wire[6:0] T13;
  wire[6:0] T14;
  wire[21:0] T15;
  wire[21:0] T50;
  wire T16;
  wire[43:0] T17;
  wire[21:0] T18;
  wire[21:0] T51;
  wire T19;
  wire[21:0] T20;
  wire[21:0] T52;
  wire T21;
  wire[87:0] T22;
  wire[87:0] T23;
  wire[43:0] T24;
  wire[21:0] wdata;
  wire[21:0] T25;
  wire[1:0] T26;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T27;
  wire[19:0] T28;
  wire[19:0] rstVal_tag;
  wire[43:0] T29;
  wire T30;
  wire[5:0] T53;
  wire[6:0] waddr;
  wire[6:0] T54;
  reg [5:0] R31;
  wire[5:0] T32;
  wire[21:0] T33;
  wire[43:0] T34;
  wire[21:0] T35;
  wire[21:0] T36;
  wire[19:0] T37;
  wire[1:0] T38;
  wire[19:0] T39;
  wire[1:0] T40;
  wire[19:0] T41;
  wire[1:0] T42;
  wire[19:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    rst_cnt = {1{$random}};
    R31 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = tags[1'h1:1'h0];
  assign tags = T1;
  assign T1 = {T34, T2};
  assign T2 = {T33, T3};
  assign T3 = T4[5'h15:1'h0];
  MetadataArray_tag_arr tag_arr (
    .CLK(clk),
    .W0A(T53),
    .W0E(T30),
    .W0I(T22),
    .W0M(T6),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(T4)
  );
  assign T6 = T7;
  assign T7 = {T17, T8};
  assign T8 = {T15, T9};
  assign T9 = 22'h0 - T48;
  assign T48 = {21'h0, T10};
  assign T10 = T11[1'h0:1'h0];
  assign T11 = rst ? 4'hf : T12;
  assign T12 = io_write_bits_way_en;
  assign rst = rst_cnt < 7'h40;
  assign T49 = reset ? 7'h0 : T13;
  assign T13 = rst ? T14 : rst_cnt;
  assign T14 = rst_cnt + 7'h1;
  assign T15 = 22'h0 - T50;
  assign T50 = {21'h0, T16};
  assign T16 = T11[1'h1:1'h1];
  assign T17 = {T20, T18};
  assign T18 = 22'h0 - T51;
  assign T51 = {21'h0, T19};
  assign T19 = T11[2'h2:2'h2];
  assign T20 = 22'h0 - T52;
  assign T52 = {21'h0, T21};
  assign T21 = T11[2'h3:2'h3];
  assign T22 = T23;
  assign T23 = {T29, T24};
  assign T24 = {wdata, wdata};
  assign wdata = T25;
  assign T25 = {T28, T26};
  assign T26 = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign rstVal_coh_state = T27;
  assign T27 = 2'h0;
  assign T28 = rst ? rstVal_tag : io_write_bits_data_tag;
  assign rstVal_tag = 20'h0;
  assign T29 = {wdata, wdata};
  assign T30 = rst | io_write_valid;
  assign T53 = waddr[3'h5:1'h0];
  assign waddr = rst ? rst_cnt : T54;
  assign T54 = {1'h0, io_write_bits_idx};
  assign T32 = io_read_valid ? io_read_bits_idx : R31;
  assign T33 = T4[6'h2b:5'h16];
  assign T34 = {T36, T35};
  assign T35 = T4[7'h41:6'h2c];
  assign T36 = T4[7'h57:7'h42];
  assign io_resp_0_tag = T37;
  assign T37 = tags[5'h15:2'h2];
  assign io_resp_1_coh_state = T38;
  assign T38 = tags[5'h17:5'h16];
  assign io_resp_1_tag = T39;
  assign T39 = tags[6'h2b:5'h18];
  assign io_resp_2_coh_state = T40;
  assign T40 = tags[6'h2d:6'h2c];
  assign io_resp_2_tag = T41;
  assign T41 = tags[7'h41:6'h2e];
  assign io_resp_3_coh_state = T42;
  assign T42 = tags[7'h43:7'h42];
  assign io_resp_3_tag = T43;
  assign T43 = tags[7'h57:7'h44];
  assign io_write_ready = T44;
  assign T44 = rst ^ 1'h1;
  assign io_read_ready = T45;
  assign T45 = T47 & T46;
  assign T46 = io_write_valid ^ 1'h1;
  assign T47 = rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else if(rst) begin
      rst_cnt <= T14;
    end
    if(io_read_valid) begin
      R31 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_0(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [5:0] io_in_4_bits_idx,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [5:0] io_in_3_bits_idx,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [5:0] io_in_2_bits_idx,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[5:0] T3;
  wire[5:0] T4;
  wire[5:0] T5;
  wire T6;
  wire[2:0] T7;
  wire[5:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 3'h0 : T0;
  assign T0 = io_in_1_valid ? 3'h1 : T1;
  assign T1 = io_in_2_valid ? 3'h2 : T2;
  assign T2 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_idx = T3;
  assign T3 = T11 ? io_in_4_bits_idx : T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = chosen;
  assign T8 = T9 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T9 = T7[1'h0:1'h0];
  assign T10 = T7[1'h1:1'h1];
  assign T11 = T7[2'h2:2'h2];
  assign io_out_valid = T12;
  assign T12 = T19 ? io_in_4_valid : T13;
  assign T13 = T18 ? T16 : T14;
  assign T14 = T15 ? io_in_1_valid : io_in_0_valid;
  assign T15 = T7[1'h0:1'h0];
  assign T16 = T17 ? io_in_3_valid : io_in_2_valid;
  assign T17 = T7[1'h0:1'h0];
  assign T18 = T7[1'h1:1'h1];
  assign T19 = T7[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T25;
  assign T25 = T26 & io_out_ready;
  assign T26 = T27 ^ 1'h1;
  assign T27 = T28 | io_in_2_valid;
  assign T28 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T29;
  assign T29 = T30 & io_out_ready;
  assign T30 = T31 ^ 1'h1;
  assign T31 = T32 | io_in_3_valid;
  assign T32 = T33 | io_in_2_valid;
  assign T33 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input [3:0] io_read_bits_way_en,
    input [11:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input [3:0] io_write_bits_way_en,
    input [11:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [127:0] io_write_bits_data,
    output[127:0] io_resp_3,
    output[127:0] io_resp_2,
    output[127:0] io_resp_1,
    output[127:0] io_resp_0
);

  wire[127:0] T0;
  wire[127:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[127:0] T4;
  wire[127:0] T5;
  wire[127:0] T6;
  wire[63:0] T7;
  wire[127:0] T8;
  wire T28;
  wire T29;
  wire[1:0] T30;
  wire[7:0] raddr;
  wire[127:0] T10;
  wire[127:0] T11;
  wire[127:0] T12;
  wire[63:0] T13;
  wire[63:0] T140;
  wire T14;
  wire[1:0] T15;
  wire[63:0] T16;
  wire[63:0] T141;
  wire T17;
  wire[127:0] T18;
  wire[127:0] T19;
  wire[63:0] T20;
  wire[63:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[7:0] waddr;
  reg [7:0] R26;
  wire[7:0] T27;
  wire[63:0] T31;
  wire T32;
  wire T33;
  reg [11:0] R34;
  wire[11:0] T35;
  wire[63:0] T36;
  wire[127:0] T37;
  wire[127:0] T38;
  wire[127:0] T39;
  wire[63:0] T40;
  wire[127:0] T41;
  wire T60;
  wire T61;
  wire[127:0] T43;
  wire[127:0] T44;
  wire[127:0] T45;
  wire[63:0] T46;
  wire[63:0] T142;
  wire T47;
  wire[63:0] T48;
  wire[63:0] T143;
  wire T49;
  wire[127:0] T50;
  wire[127:0] T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  reg [7:0] R58;
  wire[7:0] T59;
  wire[63:0] T62;
  wire[127:0] T63;
  wire[127:0] T64;
  wire[63:0] T65;
  wire[63:0] T66;
  wire T67;
  wire T68;
  wire[63:0] T69;
  wire[127:0] T70;
  wire[127:0] T71;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[127:0] T74;
  wire[127:0] T75;
  wire[127:0] T76;
  wire[63:0] T77;
  wire[127:0] T78;
  wire T98;
  wire T99;
  wire[1:0] T100;
  wire[127:0] T80;
  wire[127:0] T81;
  wire[127:0] T82;
  wire[63:0] T83;
  wire[63:0] T144;
  wire T84;
  wire[1:0] T85;
  wire[63:0] T86;
  wire[63:0] T145;
  wire T87;
  wire[127:0] T88;
  wire[127:0] T89;
  wire[63:0] T90;
  wire[63:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  reg [7:0] R96;
  wire[7:0] T97;
  wire[63:0] T101;
  wire T102;
  wire T103;
  reg [11:0] R104;
  wire[11:0] T105;
  wire[63:0] T106;
  wire[127:0] T107;
  wire[127:0] T108;
  wire[127:0] T109;
  wire[63:0] T110;
  wire[127:0] T111;
  wire T130;
  wire T131;
  wire[127:0] T113;
  wire[127:0] T114;
  wire[127:0] T115;
  wire[63:0] T116;
  wire[63:0] T146;
  wire T117;
  wire[63:0] T118;
  wire[63:0] T147;
  wire T119;
  wire[127:0] T120;
  wire[127:0] T121;
  wire[63:0] T122;
  wire[63:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  reg [7:0] R128;
  wire[7:0] T129;
  wire[63:0] T132;
  wire[127:0] T133;
  wire[127:0] T134;
  wire[63:0] T135;
  wire[63:0] T136;
  wire T137;
  wire T138;
  wire[63:0] T139;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R26 = {1{$random}};
    R34 = {1{$random}};
    R58 = {1{$random}};
    R96 = {1{$random}};
    R104 = {1{$random}};
    R128 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0 = T0;
  assign T0 = T1;
  assign T1 = {T36, T2};
  assign T2 = T32 ? T36 : T3;
  assign T3 = T4[6'h3f:1'h0];
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = {T31, T7};
  assign T7 = T8[6'h3f:1'h0];
  assign T28 = T29 & io_read_valid;
  assign T29 = T30 != 2'h0;
  assign T30 = io_read_bits_way_en[1'h1:1'h0];
  assign raddr = io_read_bits_addr >> 3'h4;
  DataArray_T9 T9 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T22),
    .W0I(T18),
    .W0M(T11),
    .R1A(raddr),
    .R1E(T28),
    .R1O(T8)
  );
  assign T11 = T12;
  assign T12 = {T16, T13};
  assign T13 = 64'h0 - T140;
  assign T140 = {63'h0, T14};
  assign T14 = T15[1'h0:1'h0];
  assign T15 = io_write_bits_way_en[1'h1:1'h0];
  assign T16 = 64'h0 - T141;
  assign T141 = {63'h0, T17};
  assign T17 = T15[1'h1:1'h1];
  assign T18 = T19;
  assign T19 = {T21, T20};
  assign T20 = io_write_bits_data[6'h3f:1'h0];
  assign T21 = io_write_bits_data[6'h3f:1'h0];
  assign T22 = T24 & T23;
  assign T23 = io_write_bits_wmask[1'h0:1'h0];
  assign T24 = T25 & io_write_valid;
  assign T25 = T15 != 2'h0;
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T27 = T28 ? raddr : R26;
  assign T31 = T8[7'h7f:7'h40];
  assign T32 = T33;
  assign T33 = R34[2'h3:2'h3];
  assign T35 = io_read_valid ? io_read_bits_addr : R34;
  assign T36 = T37[6'h3f:1'h0];
  assign T37 = T38;
  assign T38 = T39;
  assign T39 = {T62, T40};
  assign T40 = T41[6'h3f:1'h0];
  assign T60 = T61 & io_read_valid;
  assign T61 = T30 != 2'h0;
  DataArray_T9 T42 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T54),
    .W0I(T50),
    .W0M(T44),
    .R1A(raddr),
    .R1E(T60),
    .R1O(T41)
  );
  assign T44 = T45;
  assign T45 = {T48, T46};
  assign T46 = 64'h0 - T142;
  assign T142 = {63'h0, T47};
  assign T47 = T15[1'h0:1'h0];
  assign T48 = 64'h0 - T143;
  assign T143 = {63'h0, T49};
  assign T49 = T15[1'h1:1'h1];
  assign T50 = T51;
  assign T51 = {T53, T52};
  assign T52 = io_write_bits_data[7'h7f:7'h40];
  assign T53 = io_write_bits_data[7'h7f:7'h40];
  assign T54 = T56 & T55;
  assign T55 = io_write_bits_wmask[1'h1:1'h1];
  assign T56 = T57 & io_write_valid;
  assign T57 = T15 != 2'h0;
  assign T59 = T60 ? raddr : R58;
  assign T62 = T41[7'h7f:7'h40];
  assign io_resp_1 = T63;
  assign T63 = T64;
  assign T64 = {T69, T65};
  assign T65 = T67 ? T69 : T66;
  assign T66 = T4[7'h7f:7'h40];
  assign T67 = T68;
  assign T68 = R34[2'h3:2'h3];
  assign T69 = T37[7'h7f:7'h40];
  assign io_resp_2 = T70;
  assign T70 = T71;
  assign T71 = {T106, T72};
  assign T72 = T102 ? T106 : T73;
  assign T73 = T74[6'h3f:1'h0];
  assign T74 = T75;
  assign T75 = T76;
  assign T76 = {T101, T77};
  assign T77 = T78[6'h3f:1'h0];
  assign T98 = T99 & io_read_valid;
  assign T99 = T100 != 2'h0;
  assign T100 = io_read_bits_way_en[2'h3:2'h2];
  DataArray_T9 T79 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T92),
    .W0I(T88),
    .W0M(T81),
    .R1A(raddr),
    .R1E(T98),
    .R1O(T78)
  );
  assign T81 = T82;
  assign T82 = {T86, T83};
  assign T83 = 64'h0 - T144;
  assign T144 = {63'h0, T84};
  assign T84 = T85[1'h0:1'h0];
  assign T85 = io_write_bits_way_en[2'h3:2'h2];
  assign T86 = 64'h0 - T145;
  assign T145 = {63'h0, T87};
  assign T87 = T85[1'h1:1'h1];
  assign T88 = T89;
  assign T89 = {T91, T90};
  assign T90 = io_write_bits_data[6'h3f:1'h0];
  assign T91 = io_write_bits_data[6'h3f:1'h0];
  assign T92 = T94 & T93;
  assign T93 = io_write_bits_wmask[1'h0:1'h0];
  assign T94 = T95 & io_write_valid;
  assign T95 = T85 != 2'h0;
  assign T97 = T98 ? raddr : R96;
  assign T101 = T78[7'h7f:7'h40];
  assign T102 = T103;
  assign T103 = R104[2'h3:2'h3];
  assign T105 = io_read_valid ? io_read_bits_addr : R104;
  assign T106 = T107[6'h3f:1'h0];
  assign T107 = T108;
  assign T108 = T109;
  assign T109 = {T132, T110};
  assign T110 = T111[6'h3f:1'h0];
  assign T130 = T131 & io_read_valid;
  assign T131 = T100 != 2'h0;
  DataArray_T9 T112 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T124),
    .W0I(T120),
    .W0M(T114),
    .R1A(raddr),
    .R1E(T130),
    .R1O(T111)
  );
  assign T114 = T115;
  assign T115 = {T118, T116};
  assign T116 = 64'h0 - T146;
  assign T146 = {63'h0, T117};
  assign T117 = T85[1'h0:1'h0];
  assign T118 = 64'h0 - T147;
  assign T147 = {63'h0, T119};
  assign T119 = T85[1'h1:1'h1];
  assign T120 = T121;
  assign T121 = {T123, T122};
  assign T122 = io_write_bits_data[7'h7f:7'h40];
  assign T123 = io_write_bits_data[7'h7f:7'h40];
  assign T124 = T126 & T125;
  assign T125 = io_write_bits_wmask[1'h1:1'h1];
  assign T126 = T127 & io_write_valid;
  assign T127 = T85 != 2'h0;
  assign T129 = T130 ? raddr : R128;
  assign T132 = T111[7'h7f:7'h40];
  assign io_resp_3 = T133;
  assign T133 = T134;
  assign T134 = {T139, T135};
  assign T135 = T137 ? T139 : T136;
  assign T136 = T74[7'h7f:7'h40];
  assign T137 = T138;
  assign T138 = R104[2'h3:2'h3];
  assign T139 = T107[7'h7f:7'h40];
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T28) begin
      R26 <= raddr;
    end
    if(io_read_valid) begin
      R34 <= io_read_bits_addr;
    end
    if(T60) begin
      R58 <= raddr;
    end
    if(T98) begin
      R96 <= raddr;
    end
    if(io_read_valid) begin
      R104 <= io_read_bits_addr;
    end
    if(T130) begin
      R128 <= raddr;
    end
  end
endmodule

module Arbiter_2(
    output io_in_3_ready,
    input  io_in_3_valid,
    input [3:0] io_in_3_bits_way_en,
    input [11:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [3:0] io_in_2_bits_way_en,
    input [11:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[11:0] T2;
  wire[11:0] T3;
  wire T4;
  wire[1:0] T5;
  wire[11:0] T6;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire T11;
  wire[3:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 2'h0 : T0;
  assign T0 = io_in_1_valid ? 2'h1 : T1;
  assign T1 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T2;
  assign T2 = T8 ? T6 : T3;
  assign T3 = T4 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T4 = T5[1'h0:1'h0];
  assign T5 = chosen;
  assign T6 = T7 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T7 = T5[1'h0:1'h0];
  assign T8 = T5[1'h1:1'h1];
  assign io_out_bits_way_en = T9;
  assign T9 = T14 ? T12 : T10;
  assign T10 = T11 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T11 = T5[1'h0:1'h0];
  assign T12 = T13 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T13 = T5[1'h0:1'h0];
  assign T14 = T5[1'h1:1'h1];
  assign io_out_valid = T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T5[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T5[1'h0:1'h0];
  assign T20 = T5[1'h1:1'h1];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T21;
  assign T21 = T22 & io_out_ready;
  assign T22 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = T25 ^ 1'h1;
  assign T25 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T28 ^ 1'h1;
  assign T28 = T29 | io_in_2_valid;
  assign T29 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[127:0] T0;
  wire T1;
  wire[1:0] T2;
  wire[11:0] T3;
  wire[3:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T0;
  assign T0 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T1 = chosen;
  assign io_out_bits_wmask = T2;
  assign T2 = T1 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T3;
  assign T3 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T4;
  assign T4 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [4:0] io_cmd,
    input [2:0] io_typ,
    input [63:0] io_lhs,
    input [63:0] io_rhs,
    output[63:0] io_out
);

  wire[63:0] T121;
  wire[87:0] T0;
  wire[87:0] T1;
  wire[87:0] T122;
  wire[87:0] T2;
  wire[87:0] wmask;
  wire[87:0] T3;
  wire[47:0] T4;
  wire[23:0] T5;
  wire[15:0] T6;
  wire[7:0] T7;
  wire[7:0] T123;
  wire T8;
  wire[10:0] T9;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[10:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[10:0] T124;
  wire[8:0] T18;
  wire[2:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[10:0] T125;
  wire[7:0] T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T126;
  wire T30;
  wire[7:0] T31;
  wire[7:0] T127;
  wire T32;
  wire[23:0] T33;
  wire[15:0] T34;
  wire[7:0] T35;
  wire[7:0] T128;
  wire T36;
  wire[7:0] T37;
  wire[7:0] T129;
  wire T38;
  wire[7:0] T39;
  wire[7:0] T130;
  wire T40;
  wire[39:0] T41;
  wire[23:0] T42;
  wire[15:0] T43;
  wire[7:0] T44;
  wire[7:0] T131;
  wire T45;
  wire[7:0] T46;
  wire[7:0] T132;
  wire T47;
  wire[7:0] T48;
  wire[7:0] T133;
  wire T49;
  wire[15:0] T50;
  wire[7:0] T51;
  wire[7:0] T134;
  wire T52;
  wire[7:0] T53;
  wire[7:0] T135;
  wire T54;
  wire[87:0] T55;
  wire[87:0] T136;
  wire[63:0] out;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  wire[63:0] T60;
  wire[63:0] T61;
  wire[63:0] T62;
  wire[63:0] T63;
  wire[31:0] T64;
  wire[63:0] T65;
  wire[31:0] T66;
  wire[15:0] T67;
  wire[63:0] T68;
  wire[31:0] T69;
  wire[15:0] T70;
  wire[7:0] T71;
  wire T72;
  wire max;
  wire T73;
  wire T74;
  wire min;
  wire T75;
  wire T76;
  wire less;
  wire T77;
  wire cmp_rhs;
  wire T78;
  wire[63:0] rhs;
  wire[63:0] T79;
  wire[31:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire word;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire cmp_lhs;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire sgned;
  wire T96;
  wire T97;
  wire lt;
  wire T98;
  wire T99;
  wire lt_lo;
  wire[31:0] T100;
  wire[31:0] T101;
  wire eq_hi;
  wire[31:0] T102;
  wire[31:0] T103;
  wire lt_hi;
  wire[31:0] T104;
  wire[31:0] T105;
  wire T106;
  wire T107;
  wire T108;
  wire[63:0] T109;
  wire T110;
  wire[63:0] T111;
  wire T112;
  wire[63:0] T113;
  wire T114;
  wire[63:0] adder_out;
  wire[63:0] T115;
  wire[63:0] mask;
  wire[63:0] T137;
  wire[31:0] T116;
  wire T117;
  wire[63:0] T118;
  wire[63:0] T119;
  wire T120;


  assign io_out = T121;
  assign T121 = T0[6'h3f:1'h0];
  assign T0 = T55 | T1;
  assign T1 = T2 & T122;
  assign T122 = {24'h0, io_lhs};
  assign T2 = ~ wmask;
  assign wmask = T3;
  assign T3 = {T41, T4};
  assign T4 = {T33, T5};
  assign T5 = {T31, T6};
  assign T6 = {T29, T7};
  assign T7 = 8'h0 - T123;
  assign T123 = {7'h0, T8};
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T26 ? T125 : T10;
  assign T10 = T21 ? T124 : T11;
  assign T11 = T15 ? T12 : 11'hff;
  assign T12 = 4'hf << T13;
  assign T13 = {T14, 2'h0};
  assign T14 = io_addr[2'h2:2'h2];
  assign T15 = T17 | T16;
  assign T16 = io_typ == 3'h6;
  assign T17 = io_typ == 3'h2;
  assign T124 = {2'h0, T18};
  assign T18 = 2'h3 << T19;
  assign T19 = {T20, 1'h0};
  assign T20 = io_addr[2'h2:1'h1];
  assign T21 = T23 | T22;
  assign T22 = io_typ == 3'h5;
  assign T23 = io_typ == 3'h1;
  assign T125 = {3'h0, T24};
  assign T24 = 1'h1 << T25;
  assign T25 = io_addr[2'h2:1'h0];
  assign T26 = T28 | T27;
  assign T27 = io_typ == 3'h4;
  assign T28 = io_typ == 3'h0;
  assign T29 = 8'h0 - T126;
  assign T126 = {7'h0, T30};
  assign T30 = T9[1'h1:1'h1];
  assign T31 = 8'h0 - T127;
  assign T127 = {7'h0, T32};
  assign T32 = T9[2'h2:2'h2];
  assign T33 = {T39, T34};
  assign T34 = {T37, T35};
  assign T35 = 8'h0 - T128;
  assign T128 = {7'h0, T36};
  assign T36 = T9[2'h3:2'h3];
  assign T37 = 8'h0 - T129;
  assign T129 = {7'h0, T38};
  assign T38 = T9[3'h4:3'h4];
  assign T39 = 8'h0 - T130;
  assign T130 = {7'h0, T40};
  assign T40 = T9[3'h5:3'h5];
  assign T41 = {T50, T42};
  assign T42 = {T48, T43};
  assign T43 = {T46, T44};
  assign T44 = 8'h0 - T131;
  assign T131 = {7'h0, T45};
  assign T45 = T9[3'h6:3'h6];
  assign T46 = 8'h0 - T132;
  assign T132 = {7'h0, T47};
  assign T47 = T9[3'h7:3'h7];
  assign T48 = 8'h0 - T133;
  assign T133 = {7'h0, T49};
  assign T49 = T9[4'h8:4'h8];
  assign T50 = {T53, T51};
  assign T51 = 8'h0 - T134;
  assign T134 = {7'h0, T52};
  assign T52 = T9[4'h9:4'h9];
  assign T53 = 8'h0 - T135;
  assign T135 = {7'h0, T54};
  assign T54 = T9[4'ha:4'ha];
  assign T55 = wmask & T136;
  assign T136 = {24'h0, out};
  assign out = T120 ? adder_out : T56;
  assign T56 = T114 ? T113 : T57;
  assign T57 = T112 ? T111 : T58;
  assign T58 = T110 ? T109 : T59;
  assign T59 = T72 ? io_lhs : T60;
  assign T60 = T26 ? T68 : T61;
  assign T61 = T21 ? T65 : T62;
  assign T62 = T15 ? T63 : io_rhs;
  assign T63 = {T64, T64};
  assign T64 = io_rhs[5'h1f:1'h0];
  assign T65 = {T66, T66};
  assign T66 = {T67, T67};
  assign T67 = io_rhs[4'hf:1'h0];
  assign T68 = {T69, T69};
  assign T69 = {T70, T70};
  assign T70 = {T71, T71};
  assign T71 = io_rhs[3'h7:1'h0];
  assign T72 = less ? min : max;
  assign max = T74 | T73;
  assign T73 = io_cmd == 5'hf;
  assign T74 = io_cmd == 5'hd;
  assign min = T76 | T75;
  assign T75 = io_cmd == 5'he;
  assign T76 = io_cmd == 5'hc;
  assign less = T108 ? lt : T77;
  assign T77 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T82 ? T81 : T78;
  assign T78 = rhs[6'h3f:6'h3f];
  assign rhs = T15 ? T79 : io_rhs;
  assign T79 = {T80, T80};
  assign T80 = io_rhs[5'h1f:1'h0];
  assign T81 = rhs[5'h1f:5'h1f];
  assign T82 = word & T83;
  assign T83 = T84 ^ 1'h1;
  assign T84 = io_addr[2'h2:2'h2];
  assign word = T86 | T85;
  assign T85 = io_typ == 3'h4;
  assign T86 = T88 | T87;
  assign T87 = io_typ == 3'h0;
  assign T88 = T90 | T89;
  assign T89 = io_typ == 3'h6;
  assign T90 = io_typ == 3'h2;
  assign cmp_lhs = T93 ? T92 : T91;
  assign T91 = io_lhs[6'h3f:6'h3f];
  assign T92 = io_lhs[5'h1f:5'h1f];
  assign T93 = word & T94;
  assign T94 = T95 ^ 1'h1;
  assign T95 = io_addr[2'h2:2'h2];
  assign sgned = T97 | T96;
  assign T96 = io_cmd == 5'hd;
  assign T97 = io_cmd == 5'hc;
  assign lt = word ? T106 : T98;
  assign T98 = lt_hi | T99;
  assign T99 = eq_hi & lt_lo;
  assign lt_lo = T101 < T100;
  assign T100 = rhs[5'h1f:1'h0];
  assign T101 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T103 == T102;
  assign T102 = rhs[6'h3f:6'h20];
  assign T103 = io_lhs[6'h3f:6'h20];
  assign lt_hi = T105 < T104;
  assign T104 = rhs[6'h3f:6'h20];
  assign T105 = io_lhs[6'h3f:6'h20];
  assign T106 = T107 ? lt_hi : lt_lo;
  assign T107 = io_addr[2'h2:2'h2];
  assign T108 = cmp_lhs == cmp_rhs;
  assign T109 = io_lhs ^ rhs;
  assign T110 = io_cmd == 5'h9;
  assign T111 = io_lhs | rhs;
  assign T112 = io_cmd == 5'ha;
  assign T113 = io_lhs & rhs;
  assign T114 = io_cmd == 5'hb;
  assign adder_out = T118 + T115;
  assign T115 = rhs & mask;
  assign mask = 64'hffffffffffffffff ^ T137;
  assign T137 = {32'h0, T116};
  assign T116 = T117 << 5'h1f;
  assign T117 = io_addr[2'h2:2'h2];
  assign T118 = T119;
  assign T119 = io_lhs & mask;
  assign T120 = io_cmd == 5'h8;
endmodule

module LockingArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_r_type,
    input  io_in_1_bits_voluntary,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_r_type,
    input  io_in_0_bits_voluntary,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_r_type,
    output io_out_bits_voluntary,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  reg  lockIdx;
  wire T35;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  reg  locked;
  wire T36;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  reg [1:0] R18;
  wire[1:0] T37;
  wire[1:0] T19;
  wire[127:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[1:0] T24;
  wire[25:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R18 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid == 1'h0;
  assign T35 = reset ? 1'h1 : T1;
  assign T1 = T4 ? T2 : lockIdx;
  assign T2 = T3 == 1'h0;
  assign T3 = io_in_0_ready & io_in_0_valid;
  assign T4 = T6 & T5;
  assign T5 = locked ^ 1'h1;
  assign T6 = T12 & T7;
  assign T7 = T9 | T8;
  assign T8 = 3'h2 == io_out_bits_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h1 == io_out_bits_r_type;
  assign T11 = 3'h0 == io_out_bits_r_type;
  assign T12 = io_out_ready & io_out_valid;
  assign T36 = reset ? 1'h0 : T13;
  assign T13 = T15 ? 1'h0 : T14;
  assign T14 = T4 ? 1'h1 : locked;
  assign T15 = T12 & T16;
  assign T16 = T17 == 2'h0;
  assign T17 = R18 + 2'h1;
  assign T37 = reset ? 2'h0 : T19;
  assign T19 = T6 ? T17 : R18;
  assign io_out_bits_data = T20;
  assign T20 = T21 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T21 = chosen;
  assign io_out_bits_voluntary = T22;
  assign T22 = T21 ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign io_out_bits_r_type = T23;
  assign T23 = T21 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign io_out_bits_client_xact_id = T24;
  assign T24 = T21 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T25;
  assign T25 = T21 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_bits_addr_beat = T26;
  assign T26 = T21 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T27;
  assign T27 = T21 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = locked ? T30 : 1'h1;
  assign T30 = lockIdx == 1'h0;
  assign io_in_1_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = locked ? T34 : T33;
  assign T33 = io_in_0_valid ^ 1'h1;
  assign T34 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T4) begin
      lockIdx <= T2;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h0;
    end else if(T4) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T6) begin
      R18 <= T17;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input [39:0] io_cpu_req_bits_addr,
    input [8:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    input [2:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_kill,
    input  io_cpu_req_bits_phys,
    input [63:0] io_cpu_req_bits_data,
    output io_cpu_resp_valid,
    output[39:0] io_cpu_resp_bits_addr,
    output[8:0] io_cpu_resp_bits_tag,
    output[4:0] io_cpu_resp_bits_cmd,
    output[2:0] io_cpu_resp_bits_typ,
    output[63:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data_word_bypass,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[8:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_invalidate_lr,
    output io_cpu_ordered,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[1:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [25:0] io_mem_probe_bits_addr_block,
    input [1:0] io_mem_probe_bits_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[1:0] io_mem_release_bits_addr_beat,
    output[25:0] io_mem_release_bits_addr_block,
    output[1:0] io_mem_release_bits_client_xact_id,
    output[2:0] io_mem_release_bits_r_type,
    output io_mem_release_bits_voluntary,
    output[127:0] io_mem_release_bits_data
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg  R4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  reg [63:0] s2_req_data;
  wire[63:0] T17;
  wire[63:0] T18;
  wire[63:0] T19;
  reg  s1_replay;
  wire T568;
  wire T20;
  wire T21;
  wire s1_write;
  wire T22;
  wire T23;
  reg [4:0] s1_req_cmd;
  wire[4:0] T24;
  wire[4:0] T25;
  wire[4:0] T26;
  reg [4:0] s2_req_cmd;
  wire[4:0] T27;
  wire s2_recycle;
  wire T28;
  reg  s2_recycle_next;
  wire T569;
  wire T29;
  wire T30;
  reg  s1_valid;
  wire T570;
  wire T31;
  wire s2_recycle_ecc;
  wire s2_data_correctable;
  wire[1:0] T32;
  wire T33;
  wire s2_hit;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire[1:0] T47;
  reg [1:0] R48;
  wire[1:0] T49;
  wire T50;
  reg [3:0] s2_tag_match_way;
  wire[3:0] T51;
  wire[3:0] s1_tag_match_way;
  wire[3:0] T52;
  wire[1:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire[3:0] s1_tag_eq_way;
  wire[3:0] T57;
  wire[1:0] T58;
  wire T59;
  wire[19:0] T60;
  wire[31:0] s1_addr;
  wire[11:0] T61;
  reg [39:0] s1_req_addr;
  wire[39:0] T62;
  wire[39:0] T63;
  wire[39:0] T64;
  wire[39:0] T65;
  wire[39:0] T66;
  wire[39:0] T571;
  wire[31:0] T67;
  wire[25:0] T68;
  wire[39:0] T572;
  wire[31:0] T69;
  wire[25:0] T70;
  reg [39:0] s2_req_addr;
  wire[39:0] T71;
  wire[39:0] T573;
  wire T72;
  wire[19:0] T73;
  wire[1:0] T74;
  wire T75;
  wire[19:0] T76;
  wire T77;
  wire[19:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire[1:0] T89;
  wire[1:0] T90;
  wire[1:0] T91;
  reg [1:0] R92;
  wire[1:0] T93;
  wire T94;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[1:0] T97;
  reg [1:0] R98;
  wire[1:0] T99;
  wire T100;
  wire[1:0] T101;
  wire[1:0] T102;
  reg [1:0] R103;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire s2_tag_match;
  wire T127;
  wire s2_replay;
  wire T128;
  reg  R129;
  wire T574;
  reg  s2_valid;
  wire T575;
  wire s1_valid_masked;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  reg  s1_clk_en;
  reg [63:0] s1_req_data;
  wire[63:0] T135;
  wire[63:0] T136;
  wire[63:0] T137;
  wire T138;
  reg  s1_recycled;
  wire T576;
  wire T139;
  wire[63:0] T577;
  wire[127:0] s2_data_word;
  wire[127:0] s2_data_word_prebypass;
  wire[127:0] s2_data_uncorrected;
  wire[127:0] T140;
  wire[63:0] T141;
  wire[127:0] s2_data_muxed;
  wire[127:0] T142;
  wire[127:0] s2_data_3;
  wire[127:0] T143;
  wire[127:0] T144;
  reg [63:0] R145;
  wire[63:0] T578;
  wire[127:0] T146;
  wire[127:0] T579;
  wire[127:0] T147;
  wire T148;
  wire T149;
  reg [63:0] R150;
  wire[63:0] T151;
  wire[63:0] T152;
  wire T153;
  wire s1_writeback;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire[127:0] T158;
  wire[127:0] T159;
  wire[127:0] s2_data_2;
  wire[127:0] T160;
  wire[127:0] T161;
  reg [63:0] R162;
  wire[63:0] T580;
  wire[127:0] T163;
  wire[127:0] T581;
  wire[127:0] T164;
  wire T165;
  wire T166;
  reg [63:0] R167;
  wire[63:0] T168;
  wire[63:0] T169;
  wire T170;
  wire T171;
  wire[127:0] T172;
  wire[127:0] T173;
  wire[127:0] s2_data_1;
  wire[127:0] T174;
  wire[127:0] T175;
  reg [63:0] R176;
  wire[63:0] T582;
  wire[127:0] T177;
  wire[127:0] T583;
  wire[127:0] T178;
  wire T179;
  wire T180;
  reg [63:0] R181;
  wire[63:0] T182;
  wire[63:0] T183;
  wire T184;
  wire T185;
  wire[127:0] T186;
  wire[127:0] s2_data_0;
  wire[127:0] T187;
  wire[127:0] T188;
  reg [63:0] R189;
  wire[63:0] T584;
  wire[127:0] T190;
  wire[127:0] T585;
  wire[127:0] T191;
  wire T192;
  wire T193;
  reg [63:0] R194;
  wire[63:0] T195;
  wire[63:0] T196;
  wire T197;
  wire T198;
  wire[63:0] T199;
  wire[127:0] T586;
  reg [63:0] s2_store_bypass_data;
  wire[63:0] T200;
  wire[63:0] T201;
  wire[63:0] T202;
  reg [63:0] s4_req_data;
  wire[63:0] T203;
  wire T204;
  reg  s3_valid;
  wire T587;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire s2_sc_fail;
  wire T215;
  wire s2_lrsc_addr_match;
  wire T216;
  wire[33:0] T217;
  reg [33:0] lrsc_addr;
  wire[33:0] T218;
  wire[33:0] T219;
  wire T220;
  wire s2_lr;
  wire T221;
  wire T222;
  wire s2_valid_masked;
  wire T223;
  wire T224;
  wire s2_nack;
  wire s2_nack_miss;
  wire T225;
  wire T226;
  wire T227;
  wire s2_nack_victim;
  reg  s2_nack_hit;
  wire T228;
  wire s1_nack;
  wire T229;
  wire T230;
  wire T231;
  wire[5:0] T232;
  wire T233;
  wire T234;
  wire lrsc_valid;
  reg [4:0] lrsc_count;
  wire[4:0] T588;
  wire[4:0] T235;
  wire[4:0] T236;
  wire[4:0] T237;
  wire[4:0] T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire s2_sc;
  wire T243;
  wire T244;
  reg [63:0] s3_req_data;
  wire[63:0] T589;
  wire[127:0] T245;
  wire[127:0] T590;
  wire[63:0] T246;
  wire[127:0] T247;
  wire[127:0] T591;
  wire[127:0] s2_data_corrected;
  wire[127:0] T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  reg [4:0] s3_req_cmd;
  wire[4:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[36:0] T270;
  reg [39:0] s3_req_addr;
  wire[39:0] T271;
  wire[36:0] T592;
  wire[28:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire[36:0] T283;
  wire[36:0] T593;
  wire[28:0] T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  reg [4:0] s4_req_cmd;
  wire[4:0] T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[36:0] T301;
  reg [39:0] s4_req_addr;
  wire[39:0] T302;
  wire[36:0] T594;
  wire[28:0] T303;
  reg  s4_valid;
  wire T595;
  wire T304;
  reg  s2_store_bypass;
  wire T305;
  wire T306;
  reg [2:0] s2_req_typ;
  wire[2:0] T307;
  reg [2:0] s1_req_typ;
  wire[2:0] T308;
  wire[2:0] T309;
  wire[2:0] T310;
  wire[5:0] T596;
  wire[127:0] T311;
  wire[1:0] rowWMask;
  wire rowIdx;
  wire T312;
  wire[11:0] T597;
  reg [3:0] s3_way;
  wire[3:0] T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire[11:0] T598;
  wire[11:0] T599;
  wire[11:0] T600;
  wire[127:0] T326;
  wire[127:0] T327;
  wire[63:0] wdata_encoded_0;
  wire[63:0] wdata_encoded_1;
  wire[5:0] T601;
  wire[33:0] T328;
  wire[5:0] T602;
  wire[33:0] T329;
  reg  s1_req_phys;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  reg  s2_req_phys;
  wire T335;
  wire[27:0] T336;
  wire T337;
  wire T338;
  wire T339;
  wire s1_readwrite;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire s1_read;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire cache_pass;
  wire[3:0] T354;
  wire[3:0] s2_replaced_way_en;
  reg [1:0] R355;
  wire[1:0] T356;
  wire[1:0] T357;
  reg [15:0] R358;
  wire[15:0] T603;
  wire[15:0] T359;
  wire[15:0] T360;
  wire[14:0] T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire[1:0] T372;
  wire[21:0] T373;
  wire[21:0] T374;
  wire[21:0] T375;
  wire[21:0] T376;
  reg [1:0] R377;
  wire[1:0] T378;
  wire T379;
  wire T380;
  wire[3:0] s1_replaced_way_en;
  wire[1:0] T381;
  reg [19:0] R382;
  wire[19:0] T383;
  wire T384;
  wire[21:0] T385;
  wire[21:0] T386;
  wire[21:0] T387;
  wire[21:0] T388;
  reg [1:0] R389;
  wire[1:0] T390;
  wire T391;
  wire T392;
  reg [19:0] R393;
  wire[19:0] T394;
  wire T395;
  wire[21:0] T396;
  wire[21:0] T397;
  wire[21:0] T398;
  wire[21:0] T399;
  reg [1:0] R400;
  wire[1:0] T401;
  wire T402;
  wire T403;
  reg [19:0] R404;
  wire[19:0] T405;
  wire T406;
  wire[21:0] T407;
  wire[21:0] T408;
  wire[21:0] T409;
  reg [1:0] R410;
  wire[1:0] T411;
  wire T412;
  wire T413;
  reg [19:0] R414;
  wire[19:0] T415;
  wire T416;
  wire[1:0] T417;
  wire[19:0] T418;
  wire[19:0] T419;
  wire[19:0] T420;
  reg  s2_req_kill;
  wire T421;
  reg  s1_req_kill;
  wire T422;
  wire T423;
  wire T424;
  reg [8:0] s2_req_tag;
  wire[8:0] T425;
  reg [8:0] s1_req_tag;
  wire[8:0] T426;
  wire[8:0] T427;
  wire[8:0] T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire misaligned;
  wire T465;
  wire T466;
  wire[2:0] T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire[1:0] T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[63:0] T484;
  wire[63:0] uncache_resp_bits_store_data;
  wire[63:0] cache_resp_bits_store_data;
  wire[63:0] T485;
  wire[31:0] T486;
  wire[31:0] T487;
  wire[31:0] T488;
  wire T489;
  wire[31:0] T490;
  wire[31:0] T491;
  wire[31:0] T492;
  wire[31:0] T604;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire uncache_resp_bits_has_data;
  wire cache_resp_bits_has_data;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire uncache_resp_bits_replay;
  wire cache_resp_bits_replay;
  wire T516;
  wire uncache_resp_bits_nack;
  wire cache_resp_bits_nack;
  wire T517;
  wire[63:0] T518;
  wire[63:0] uncache_resp_bits_data;
  wire[63:0] cache_resp_bits_data;
  wire[63:0] T519;
  wire[63:0] T605;
  wire[63:0] T520;
  wire[7:0] T521;
  wire[7:0] T522;
  wire[7:0] T523;
  wire[63:0] T524;
  wire[15:0] T525;
  wire[15:0] T526;
  wire[15:0] T527;
  wire T528;
  wire[47:0] T529;
  wire[47:0] T530;
  wire[47:0] T531;
  wire[47:0] T606;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire[7:0] T537;
  wire T538;
  wire[55:0] T539;
  wire[55:0] T540;
  wire[55:0] T541;
  wire[55:0] T607;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[2:0] T548;
  wire[2:0] uncache_resp_bits_typ;
  wire[2:0] cache_resp_bits_typ;
  wire[4:0] T549;
  wire[4:0] uncache_resp_bits_cmd;
  wire[4:0] cache_resp_bits_cmd;
  wire[8:0] T550;
  wire[8:0] uncache_resp_bits_tag;
  wire[8:0] cache_resp_bits_tag;
  wire[39:0] T551;
  wire[39:0] uncache_resp_bits_addr;
  wire[39:0] cache_resp_bits_addr;
  wire T552;
  wire uncache_resp_valid;
  wire cache_resp_valid;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  reg  block_miss;
  wire T608;
  wire T566;
  wire T567;
  wire wb_io_req_ready;
  wire wb_io_meta_read_valid;
  wire[5:0] wb_io_meta_read_bits_idx;
  wire[19:0] wb_io_meta_read_bits_tag;
  wire wb_io_data_req_valid;
  wire[3:0] wb_io_data_req_bits_way_en;
  wire[11:0] wb_io_data_req_bits_addr;
  wire wb_io_release_valid;
  wire[1:0] wb_io_release_bits_addr_beat;
  wire[25:0] wb_io_release_bits_addr_block;
  wire[1:0] wb_io_release_bits_client_xact_id;
  wire[2:0] wb_io_release_bits_r_type;
  wire wb_io_release_bits_voluntary;
  wire[127:0] wb_io_release_bits_data;
  wire prober_io_req_ready;
  wire prober_io_rep_valid;
  wire[1:0] prober_io_rep_bits_addr_beat;
  wire[25:0] prober_io_rep_bits_addr_block;
  wire[1:0] prober_io_rep_bits_client_xact_id;
  wire[2:0] prober_io_rep_bits_r_type;
  wire prober_io_rep_bits_voluntary;
  wire[127:0] prober_io_rep_bits_data;
  wire prober_io_meta_read_valid;
  wire[5:0] prober_io_meta_read_bits_idx;
  wire[19:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_write_valid;
  wire[5:0] prober_io_meta_write_bits_idx;
  wire[3:0] prober_io_meta_write_bits_way_en;
  wire[19:0] prober_io_meta_write_bits_data_tag;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire prober_io_wb_req_valid;
  wire[1:0] prober_io_wb_req_bits_addr_beat;
  wire[25:0] prober_io_wb_req_bits_addr_block;
  wire[1:0] prober_io_wb_req_bits_client_xact_id;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire prober_io_wb_req_bits_voluntary;
  wire[127:0] prober_io_wb_req_bits_data;
  wire[3:0] prober_io_wb_req_bits_way_en;
  wire meta_io_read_ready;
  wire meta_io_write_ready;
  wire[19:0] meta_io_resp_3_tag;
  wire[1:0] meta_io_resp_3_coh_state;
  wire[19:0] meta_io_resp_2_tag;
  wire[1:0] meta_io_resp_2_coh_state;
  wire[19:0] meta_io_resp_1_tag;
  wire[1:0] meta_io_resp_1_coh_state;
  wire[19:0] meta_io_resp_0_tag;
  wire[1:0] meta_io_resp_0_coh_state;
  wire metaReadArb_io_in_4_ready;
  wire metaReadArb_io_in_3_ready;
  wire metaReadArb_io_in_2_ready;
  wire metaReadArb_io_in_1_ready;
  wire metaReadArb_io_out_valid;
  wire[5:0] metaReadArb_io_out_bits_idx;
  wire metaWriteArb_io_in_1_ready;
  wire metaWriteArb_io_in_0_ready;
  wire metaWriteArb_io_out_valid;
  wire[5:0] metaWriteArb_io_out_bits_idx;
  wire[3:0] metaWriteArb_io_out_bits_way_en;
  wire[19:0] metaWriteArb_io_out_bits_data_tag;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire data_io_write_ready;
  wire[127:0] data_io_resp_3;
  wire[127:0] data_io_resp_2;
  wire[127:0] data_io_resp_1;
  wire[127:0] data_io_resp_0;
  wire readArb_io_in_3_ready;
  wire readArb_io_in_2_ready;
  wire readArb_io_in_1_ready;
  wire readArb_io_out_valid;
  wire[3:0] readArb_io_out_bits_way_en;
  wire[11:0] readArb_io_out_bits_addr;
  wire writeArb_io_in_1_ready;
  wire writeArb_io_out_valid;
  wire[3:0] writeArb_io_out_bits_way_en;
  wire[11:0] writeArb_io_out_bits_addr;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[127:0] writeArb_io_out_bits_data;
  wire[63:0] amoalu_io_out;
  wire releaseArb_io_in_1_ready;
  wire releaseArb_io_in_0_ready;
  wire releaseArb_io_out_valid;
  wire[1:0] releaseArb_io_out_bits_addr_beat;
  wire[25:0] releaseArb_io_out_bits_addr_block;
  wire[1:0] releaseArb_io_out_bits_client_xact_id;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire releaseArb_io_out_bits_voluntary;
  wire[127:0] releaseArb_io_out_bits_data;
  wire FlowThroughSerializer_io_in_ready;
  wire FlowThroughSerializer_io_out_valid;
  wire[1:0] FlowThroughSerializer_io_out_bits_addr_beat;
  wire[1:0] FlowThroughSerializer_io_out_bits_client_xact_id;
  wire[3:0] FlowThroughSerializer_io_out_bits_manager_xact_id;
  wire FlowThroughSerializer_io_out_bits_is_builtin_type;
  wire[3:0] FlowThroughSerializer_io_out_bits_g_type;
  wire[127:0] FlowThroughSerializer_io_out_bits_data;
  wire wbArb_io_in_1_ready;
  wire wbArb_io_in_0_ready;
  wire wbArb_io_out_valid;
  wire[1:0] wbArb_io_out_bits_addr_beat;
  wire[25:0] wbArb_io_out_bits_addr_block;
  wire[1:0] wbArb_io_out_bits_client_xact_id;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire wbArb_io_out_bits_voluntary;
  wire[127:0] wbArb_io_out_bits_data;
  wire[3:0] wbArb_io_out_bits_way_en;
  wire dtlb_io_req_ready;
  wire dtlb_io_resp_miss;
  wire[19:0] dtlb_io_resp_ppn;
  wire dtlb_io_resp_xcpt_ld;
  wire dtlb_io_resp_xcpt_st;
  wire dtlb_io_ptw_req_valid;
  wire[26:0] dtlb_io_ptw_req_bits_addr;
  wire[1:0] dtlb_io_ptw_req_bits_prv;
  wire dtlb_io_ptw_req_bits_store;
  wire dtlb_io_ptw_req_bits_fetch;
  wire mshrs_io_req_ready;
  wire mshrs_io_resp_valid;
  wire[39:0] mshrs_io_resp_bits_addr;
  wire[8:0] mshrs_io_resp_bits_tag;
  wire[4:0] mshrs_io_resp_bits_cmd;
  wire[2:0] mshrs_io_resp_bits_typ;
  wire[63:0] mshrs_io_resp_bits_data;
  wire mshrs_io_resp_bits_nack;
  wire mshrs_io_resp_bits_replay;
  wire mshrs_io_resp_bits_has_data;
  wire[63:0] mshrs_io_resp_bits_store_data;
  wire mshrs_io_secondary_miss;
  wire mshrs_io_mem_req_valid;
  wire[25:0] mshrs_io_mem_req_bits_addr_block;
  wire[1:0] mshrs_io_mem_req_bits_client_xact_id;
  wire[1:0] mshrs_io_mem_req_bits_addr_beat;
  wire mshrs_io_mem_req_bits_is_builtin_type;
  wire[2:0] mshrs_io_mem_req_bits_a_type;
  wire[16:0] mshrs_io_mem_req_bits_union;
  wire[127:0] mshrs_io_mem_req_bits_data;
  wire[3:0] mshrs_io_refill_way_en;
  wire[11:0] mshrs_io_refill_addr;
  wire mshrs_io_meta_read_valid;
  wire[5:0] mshrs_io_meta_read_bits_idx;
  wire mshrs_io_meta_write_valid;
  wire[5:0] mshrs_io_meta_write_bits_idx;
  wire[3:0] mshrs_io_meta_write_bits_way_en;
  wire[19:0] mshrs_io_meta_write_bits_data_tag;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire mshrs_io_replay_valid;
  wire[39:0] mshrs_io_replay_bits_addr;
  wire[8:0] mshrs_io_replay_bits_tag;
  wire[4:0] mshrs_io_replay_bits_cmd;
  wire[2:0] mshrs_io_replay_bits_typ;
  wire mshrs_io_replay_bits_kill;
  wire mshrs_io_replay_bits_phys;
  wire[63:0] mshrs_io_replay_bits_data;
  wire mshrs_io_wb_req_valid;
  wire[1:0] mshrs_io_wb_req_bits_addr_beat;
  wire[25:0] mshrs_io_wb_req_bits_addr_block;
  wire[1:0] mshrs_io_wb_req_bits_client_xact_id;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire mshrs_io_wb_req_bits_voluntary;
  wire[127:0] mshrs_io_wb_req_bits_data;
  wire[3:0] mshrs_io_wb_req_bits_way_en;
  wire mshrs_io_probe_rdy;
  wire mshrs_io_fence_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {1{$random}};
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s2_recycle_next = {1{$random}};
    s1_valid = {1{$random}};
    R48 = {1{$random}};
    s2_tag_match_way = {1{$random}};
    s1_req_addr = {2{$random}};
    s2_req_addr = {2{$random}};
    R92 = {1{$random}};
    R98 = {1{$random}};
    R103 = {1{$random}};
    R129 = {1{$random}};
    s2_valid = {1{$random}};
    s1_clk_en = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R145 = {2{$random}};
    R150 = {2{$random}};
    R162 = {2{$random}};
    R167 = {2{$random}};
    R176 = {2{$random}};
    R181 = {2{$random}};
    R189 = {2{$random}};
    R194 = {2{$random}};
    s2_store_bypass_data = {2{$random}};
    s4_req_data = {2{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_data = {2{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    R355 = {1{$random}};
    R358 = {1{$random}};
    R377 = {1{$random}};
    R382 = {1{$random}};
    R389 = {1{$random}};
    R393 = {1{$random}};
    R400 = {1{$random}};
    R404 = {1{$random}};
    R410 = {1{$random}};
    R414 = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    block_miss = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = R4 & io_cpu_resp_valid;
  assign T5 = T6 | io_cpu_xcpt_pf_st;
  assign T6 = T7 | io_cpu_xcpt_pf_ld;
  assign T7 = io_cpu_xcpt_ma_ld | io_cpu_xcpt_ma_st;
  assign T8 = writeArb_io_in_1_ready | T9;
  assign T9 = T10 ^ 1'h1;
  assign T10 = FlowThroughSerializer_io_out_bits_is_builtin_type ? T14 : T11;
  assign T11 = T13 | T12;
  assign T12 = 4'h1 == FlowThroughSerializer_io_out_bits_g_type;
  assign T13 = 4'h0 == FlowThroughSerializer_io_out_bits_g_type;
  assign T14 = T16 | T15;
  assign T15 = 4'h4 == FlowThroughSerializer_io_out_bits_g_type;
  assign T16 = 4'h5 == FlowThroughSerializer_io_out_bits_g_type;
  assign T17 = T138 ? s1_req_data : T18;
  assign T18 = T21 ? T19 : s2_req_data;
  assign T19 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T568 = reset ? 1'h0 : T20;
  assign T20 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T21 = s1_clk_en & s1_write;
  assign s1_write = T132 | T22;
  assign T22 = T131 | T23;
  assign T23 = s1_req_cmd == 5'h4;
  assign T24 = s2_recycle ? s2_req_cmd : T25;
  assign T25 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T26;
  assign T26 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T27 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T28;
  assign T28 = s2_recycle_ecc | s2_recycle_next;
  assign T569 = reset ? 1'h0 : T29;
  assign T29 = T30 ? s2_recycle_ecc : s2_recycle_next;
  assign T30 = s1_valid | s1_replay;
  assign T570 = reset ? 1'h0 : T31;
  assign T31 = io_cpu_req_ready & io_cpu_req_valid;
  assign s2_recycle_ecc = T33 & s2_data_correctable;
  assign s2_data_correctable = T32[1'h0:1'h0];
  assign T32 = 2'h0;
  assign T33 = T127 & s2_hit;
  assign s2_hit = T106 & T34;
  assign T34 = T44 == T35;
  assign T35 = T36;
  assign T36 = T37 ? 2'h3 : T44;
  assign T37 = T41 | T38;
  assign T38 = T40 | T39;
  assign T39 = s2_req_cmd == 5'h4;
  assign T40 = s2_req_cmd[2'h3:2'h3];
  assign T41 = T43 | T42;
  assign T42 = s2_req_cmd == 5'h7;
  assign T43 = s2_req_cmd == 5'h1;
  assign T44 = T45[1'h1:1'h0];
  assign T45 = T89 | T46;
  assign T46 = T50 ? T47 : 2'h0;
  assign T47 = R48;
  assign T49 = s1_clk_en ? meta_io_resp_3_coh_state : R48;
  assign T50 = s2_tag_match_way[2'h3:2'h3];
  assign T51 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T52;
  assign T52 = {T82, T53};
  assign T53 = {T79, T54};
  assign T54 = T56 & T55;
  assign T55 = meta_io_resp_0_coh_state != 2'h0;
  assign T56 = s1_tag_eq_way[1'h0:1'h0];
  assign s1_tag_eq_way = T57;
  assign T57 = {T74, T58};
  assign T58 = {T72, T59};
  assign T59 = meta_io_resp_0_tag == T60;
  assign T60 = s1_addr >> 4'hc;
  assign s1_addr = {dtlb_io_resp_ppn, T61};
  assign T61 = s1_req_addr[4'hb:1'h0];
  assign T62 = s2_recycle ? s2_req_addr : T63;
  assign T63 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T64;
  assign T64 = prober_io_meta_read_valid ? T572 : T65;
  assign T65 = wb_io_meta_read_valid ? T571 : T66;
  assign T66 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T571 = {8'h0, T67};
  assign T67 = T68 << 3'h6;
  assign T68 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T572 = {8'h0, T69};
  assign T69 = T70 << 3'h6;
  assign T70 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T71 = s1_clk_en ? T573 : s2_req_addr;
  assign T573 = {8'h0, s1_addr};
  assign T72 = meta_io_resp_1_tag == T73;
  assign T73 = s1_addr >> 4'hc;
  assign T74 = {T77, T75};
  assign T75 = meta_io_resp_2_tag == T76;
  assign T76 = s1_addr >> 4'hc;
  assign T77 = meta_io_resp_3_tag == T78;
  assign T78 = s1_addr >> 4'hc;
  assign T79 = T81 & T80;
  assign T80 = meta_io_resp_1_coh_state != 2'h0;
  assign T81 = s1_tag_eq_way[1'h1:1'h1];
  assign T82 = {T86, T83};
  assign T83 = T85 & T84;
  assign T84 = meta_io_resp_2_coh_state != 2'h0;
  assign T85 = s1_tag_eq_way[2'h2:2'h2];
  assign T86 = T88 & T87;
  assign T87 = meta_io_resp_3_coh_state != 2'h0;
  assign T88 = s1_tag_eq_way[2'h3:2'h3];
  assign T89 = T95 | T90;
  assign T90 = T94 ? T91 : 2'h0;
  assign T91 = R92;
  assign T93 = s1_clk_en ? meta_io_resp_2_coh_state : R92;
  assign T94 = s2_tag_match_way[2'h2:2'h2];
  assign T95 = T101 | T96;
  assign T96 = T100 ? T97 : 2'h0;
  assign T97 = R98;
  assign T99 = s1_clk_en ? meta_io_resp_1_coh_state : R98;
  assign T100 = s2_tag_match_way[1'h1:1'h1];
  assign T101 = T105 ? T102 : 2'h0;
  assign T102 = R103;
  assign T104 = s1_clk_en ? meta_io_resp_0_coh_state : R103;
  assign T105 = s2_tag_match_way[1'h0:1'h0];
  assign T106 = s2_tag_match & T107;
  assign T107 = T116 ? T113 : T108;
  assign T108 = T110 | T109;
  assign T109 = 2'h3 == T44;
  assign T110 = T112 | T111;
  assign T111 = 2'h2 == T44;
  assign T112 = 2'h1 == T44;
  assign T113 = T115 | T114;
  assign T114 = 2'h3 == T44;
  assign T115 = 2'h2 == T44;
  assign T116 = T118 | T117;
  assign T117 = s2_req_cmd == 5'h6;
  assign T118 = T120 | T119;
  assign T119 = s2_req_cmd == 5'h3;
  assign T120 = T124 | T121;
  assign T121 = T123 | T122;
  assign T122 = s2_req_cmd == 5'h4;
  assign T123 = s2_req_cmd[2'h3:2'h3];
  assign T124 = T126 | T125;
  assign T125 = s2_req_cmd == 5'h7;
  assign T126 = s2_req_cmd == 5'h1;
  assign s2_tag_match = s2_tag_match_way != 4'h0;
  assign T127 = s2_valid | s2_replay;
  assign s2_replay = R129 & T128;
  assign T128 = s2_req_cmd != 5'h5;
  assign T574 = reset ? 1'h0 : s1_replay;
  assign T575 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T130;
  assign T130 = io_cpu_req_bits_kill ^ 1'h1;
  assign T131 = s1_req_cmd[2'h3:2'h3];
  assign T132 = T134 | T133;
  assign T133 = s1_req_cmd == 5'h7;
  assign T134 = s1_req_cmd == 5'h1;
  assign T135 = s2_recycle ? s2_req_data : T136;
  assign T136 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T137;
  assign T137 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T138 = s1_clk_en & s1_recycled;
  assign T576 = reset ? 1'h0 : T139;
  assign T139 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T577 = s2_data_word[6'h3f:1'h0];
  assign s2_data_word = s2_store_bypass ? T586 : s2_data_word_prebypass;
  assign s2_data_word_prebypass = s2_data_uncorrected >> 7'h0;
  assign s2_data_uncorrected = T140;
  assign T140 = {T199, T141};
  assign T141 = s2_data_muxed[6'h3f:1'h0];
  assign s2_data_muxed = T158 | T142;
  assign T142 = T157 ? s2_data_3 : 128'h0;
  assign s2_data_3 = T143;
  assign T143 = T144;
  assign T144 = {R150, R145};
  assign T578 = T146[6'h3f:1'h0];
  assign T146 = T148 ? T147 : T579;
  assign T579 = {64'h0, R145};
  assign T147 = data_io_resp_3 >> 1'h0;
  assign T148 = s1_clk_en & T149;
  assign T149 = s1_tag_eq_way[2'h3:2'h3];
  assign T151 = T153 ? T152 : R150;
  assign T152 = data_io_resp_3 >> 7'h40;
  assign T153 = T148 & s1_writeback;
  assign s1_writeback = T155 & T154;
  assign T154 = s1_replay ^ 1'h1;
  assign T155 = s1_clk_en & T156;
  assign T156 = s1_valid ^ 1'h1;
  assign T157 = s2_tag_match_way[2'h3:2'h3];
  assign T158 = T172 | T159;
  assign T159 = T171 ? s2_data_2 : 128'h0;
  assign s2_data_2 = T160;
  assign T160 = T161;
  assign T161 = {R167, R162};
  assign T580 = T163[6'h3f:1'h0];
  assign T163 = T165 ? T164 : T581;
  assign T581 = {64'h0, R162};
  assign T164 = data_io_resp_2 >> 1'h0;
  assign T165 = s1_clk_en & T166;
  assign T166 = s1_tag_eq_way[2'h2:2'h2];
  assign T168 = T170 ? T169 : R167;
  assign T169 = data_io_resp_2 >> 7'h40;
  assign T170 = T165 & s1_writeback;
  assign T171 = s2_tag_match_way[2'h2:2'h2];
  assign T172 = T186 | T173;
  assign T173 = T185 ? s2_data_1 : 128'h0;
  assign s2_data_1 = T174;
  assign T174 = T175;
  assign T175 = {R181, R176};
  assign T582 = T177[6'h3f:1'h0];
  assign T177 = T179 ? T178 : T583;
  assign T583 = {64'h0, R176};
  assign T178 = data_io_resp_1 >> 1'h0;
  assign T179 = s1_clk_en & T180;
  assign T180 = s1_tag_eq_way[1'h1:1'h1];
  assign T182 = T184 ? T183 : R181;
  assign T183 = data_io_resp_1 >> 7'h40;
  assign T184 = T179 & s1_writeback;
  assign T185 = s2_tag_match_way[1'h1:1'h1];
  assign T186 = T198 ? s2_data_0 : 128'h0;
  assign s2_data_0 = T187;
  assign T187 = T188;
  assign T188 = {R194, R189};
  assign T584 = T190[6'h3f:1'h0];
  assign T190 = T192 ? T191 : T585;
  assign T585 = {64'h0, R189};
  assign T191 = data_io_resp_0 >> 1'h0;
  assign T192 = s1_clk_en & T193;
  assign T193 = s1_tag_eq_way[1'h0:1'h0];
  assign T195 = T197 ? T196 : R194;
  assign T196 = data_io_resp_0 >> 7'h40;
  assign T197 = T192 & s1_writeback;
  assign T198 = s2_tag_match_way[1'h0:1'h0];
  assign T199 = s2_data_muxed[7'h7f:7'h40];
  assign T586 = {64'h0, s2_store_bypass_data};
  assign T200 = T288 ? T201 : s2_store_bypass_data;
  assign T201 = T273 ? amoalu_io_out : T202;
  assign T202 = T259 ? s3_req_data : s4_req_data;
  assign T203 = T204 ? s3_req_data : s4_req_data;
  assign T204 = s3_valid & metaReadArb_io_out_valid;
  assign T587 = reset ? 1'h0 : T205;
  assign T205 = T213 & T206;
  assign T206 = T210 | T207;
  assign T207 = T209 | T208;
  assign T208 = s2_req_cmd == 5'h4;
  assign T209 = s2_req_cmd[2'h3:2'h3];
  assign T210 = T212 | T211;
  assign T211 = s2_req_cmd == 5'h7;
  assign T212 = s2_req_cmd == 5'h1;
  assign T213 = T243 & T214;
  assign T214 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T215;
  assign T215 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = lrsc_valid & T216;
  assign T216 = lrsc_addr == T217;
  assign T217 = s2_req_addr >> 3'h6;
  assign T218 = T220 ? T219 : lrsc_addr;
  assign T219 = s2_req_addr >> 3'h6;
  assign T220 = T221 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T221 = T222 | s2_replay;
  assign T222 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T223;
  assign T223 = s2_valid & T224;
  assign T224 = s2_nack ^ 1'h1;
  assign s2_nack = T227 | s2_nack_miss;
  assign s2_nack_miss = T226 & T225;
  assign T225 = mshrs_io_req_ready ^ 1'h1;
  assign T226 = s2_hit ^ 1'h1;
  assign T227 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T228 = T234 ? s1_nack : s2_nack_hit;
  assign s1_nack = T233 | T229;
  assign T229 = T231 & T230;
  assign T230 = prober_io_req_ready ^ 1'h1;
  assign T231 = T232 == prober_io_meta_write_bits_idx;
  assign T232 = s1_req_addr[4'hb:3'h6];
  assign T233 = T337 & dtlb_io_resp_miss;
  assign T234 = s1_valid | s1_replay;
  assign lrsc_valid = lrsc_count != 5'h0;
  assign T588 = reset ? 5'h0 : T235;
  assign T235 = io_cpu_invalidate_lr ? 5'h0 : T236;
  assign T236 = T242 ? 5'h0 : T237;
  assign T237 = T240 ? 5'h1f : T238;
  assign T238 = lrsc_valid ? T239 : lrsc_count;
  assign T239 = lrsc_count - 5'h1;
  assign T240 = T220 & T241;
  assign T241 = lrsc_valid ^ 1'h1;
  assign T242 = T221 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T243 = T244 | s2_replay;
  assign T244 = s2_valid_masked & s2_hit;
  assign T589 = T245[6'h3f:1'h0];
  assign T245 = T249 ? T247 : T590;
  assign T590 = {64'h0, T246};
  assign T246 = T249 ? s2_req_data : s3_req_data;
  assign T247 = s2_data_correctable ? s2_data_corrected : T591;
  assign T591 = {64'h0, amoalu_io_out};
  assign s2_data_corrected = T248;
  assign T248 = {T199, T141};
  assign T249 = T258 & T250;
  assign T250 = T251 | s2_data_correctable;
  assign T251 = T255 | T252;
  assign T252 = T254 | T253;
  assign T253 = s2_req_cmd == 5'h4;
  assign T254 = s2_req_cmd[2'h3:2'h3];
  assign T255 = T257 | T256;
  assign T256 = s2_req_cmd == 5'h7;
  assign T257 = s2_req_cmd == 5'h1;
  assign T258 = s2_valid | s2_replay;
  assign T259 = T268 & T260;
  assign T260 = T265 | T261;
  assign T261 = T264 | T262;
  assign T262 = s3_req_cmd == 5'h4;
  assign T263 = T249 ? s2_req_cmd : s3_req_cmd;
  assign T264 = s3_req_cmd[2'h3:2'h3];
  assign T265 = T267 | T266;
  assign T266 = s3_req_cmd == 5'h7;
  assign T267 = s3_req_cmd == 5'h1;
  assign T268 = s3_valid & T269;
  assign T269 = T592 == T270;
  assign T270 = s3_req_addr >> 2'h3;
  assign T271 = T249 ? s2_req_addr : s3_req_addr;
  assign T592 = {8'h0, T272};
  assign T272 = s1_addr >> 2'h3;
  assign T273 = T281 & T274;
  assign T274 = T278 | T275;
  assign T275 = T277 | T276;
  assign T276 = s2_req_cmd == 5'h4;
  assign T277 = s2_req_cmd[2'h3:2'h3];
  assign T278 = T280 | T279;
  assign T279 = s2_req_cmd == 5'h7;
  assign T280 = s2_req_cmd == 5'h1;
  assign T281 = T285 & T282;
  assign T282 = T593 == T283;
  assign T283 = s2_req_addr >> 2'h3;
  assign T593 = {8'h0, T284};
  assign T284 = s1_addr >> 2'h3;
  assign T285 = T287 & T286;
  assign T286 = s2_sc_fail ^ 1'h1;
  assign T287 = s2_valid_masked | s2_replay;
  assign T288 = s1_clk_en & T289;
  assign T289 = T304 | T290;
  assign T290 = T299 & T291;
  assign T291 = T296 | T292;
  assign T292 = T295 | T293;
  assign T293 = s4_req_cmd == 5'h4;
  assign T294 = T204 ? s3_req_cmd : s4_req_cmd;
  assign T295 = s4_req_cmd[2'h3:2'h3];
  assign T296 = T298 | T297;
  assign T297 = s4_req_cmd == 5'h7;
  assign T298 = s4_req_cmd == 5'h1;
  assign T299 = s4_valid & T300;
  assign T300 = T594 == T301;
  assign T301 = s4_req_addr >> 2'h3;
  assign T302 = T204 ? s3_req_addr : s4_req_addr;
  assign T594 = {8'h0, T303};
  assign T303 = s1_addr >> 2'h3;
  assign T595 = reset ? 1'h0 : s3_valid;
  assign T304 = T273 | T259;
  assign T305 = T288 ? 1'h1 : T306;
  assign T306 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T307 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T308 = s2_recycle ? s2_req_typ : T309;
  assign T309 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T310;
  assign T310 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T596 = s2_req_addr[3'h5:1'h0];
  assign T311 = {s3_req_data, s3_req_data};
  assign rowWMask = 1'h1 << rowIdx;
  assign rowIdx = T312;
  assign T312 = s3_req_addr[2'h3:2'h3];
  assign T597 = s3_req_addr[4'hb:1'h0];
  assign T313 = T249 ? s2_tag_match_way : s3_way;
  assign T314 = T316 & T315;
  assign T315 = FlowThroughSerializer_io_out_bits_client_xact_id < 2'h2;
  assign T316 = FlowThroughSerializer_io_out_valid & T317;
  assign T317 = FlowThroughSerializer_io_out_bits_is_builtin_type ? T321 : T318;
  assign T318 = T320 | T319;
  assign T319 = 4'h1 == FlowThroughSerializer_io_out_bits_g_type;
  assign T320 = 4'h0 == FlowThroughSerializer_io_out_bits_g_type;
  assign T321 = T323 | T322;
  assign T322 = 4'h4 == FlowThroughSerializer_io_out_bits_g_type;
  assign T323 = 4'h5 == FlowThroughSerializer_io_out_bits_g_type;
  assign T324 = T325 | T8;
  assign T325 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T598 = s2_req_addr[4'hb:1'h0];
  assign T599 = mshrs_io_replay_bits_addr[4'hb:1'h0];
  assign T600 = io_cpu_req_bits_addr[4'hb:1'h0];
  assign T326 = T327;
  assign T327 = {wdata_encoded_1, wdata_encoded_0};
  assign wdata_encoded_0 = writeArb_io_out_bits_data[6'h3f:1'h0];
  assign wdata_encoded_1 = writeArb_io_out_bits_data[7'h7f:7'h40];
  assign T601 = T328[3'h5:1'h0];
  assign T328 = s2_req_addr >> 3'h6;
  assign T602 = T329[3'h5:1'h0];
  assign T329 = io_cpu_req_bits_addr >> 3'h6;
  assign T330 = s2_recycle ? s2_req_phys : T331;
  assign T331 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T332;
  assign T332 = prober_io_meta_read_valid ? 1'h1 : T333;
  assign T333 = wb_io_meta_read_valid ? 1'h1 : T334;
  assign T334 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T335 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T336 = s1_req_addr >> 4'hc;
  assign T337 = T339 & T338;
  assign T338 = s1_req_phys ^ 1'h1;
  assign T339 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T343 | T340;
  assign T340 = T342 | T341;
  assign T341 = s1_req_cmd == 5'h3;
  assign T342 = s1_req_cmd == 5'h2;
  assign T343 = s1_read | s1_write;
  assign s1_read = T347 | T344;
  assign T344 = T346 | T345;
  assign T345 = s1_req_cmd == 5'h4;
  assign T346 = s1_req_cmd[2'h3:2'h3];
  assign T347 = T349 | T348;
  assign T348 = s1_req_cmd == 5'h7;
  assign T349 = T351 | T350;
  assign T350 = s1_req_cmd == 5'h6;
  assign T351 = s1_req_cmd == 5'h0;
  assign T352 = T8 & FlowThroughSerializer_io_out_valid;
  assign T353 = cache_pass ^ 1'h1;
  assign cache_pass = s2_valid | s2_replay;
  assign T354 = s2_tag_match ? s2_tag_match_way : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R355;
  assign T356 = s1_clk_en ? T357 : R355;
  assign T357 = R358[1'h1:1'h0];
  assign T603 = reset ? 16'h1 : T359;
  assign T359 = T369 ? T360 : R358;
  assign T360 = {T362, T361};
  assign T361 = R358[4'hf:1'h1];
  assign T362 = T364 ^ T363;
  assign T363 = R358[3'h5:3'h5];
  assign T364 = T366 ^ T365;
  assign T365 = R358[2'h3:2'h3];
  assign T366 = T368 ^ T367;
  assign T367 = R358[2'h2:2'h2];
  assign T368 = R358[1'h0:1'h0];
  assign T369 = T370;
  assign T370 = mshrs_io_req_ready & T429;
  assign T371 = s2_tag_match ? T417 : T372;
  assign T372 = T373[1'h1:1'h0];
  assign T373 = T385 | T374;
  assign T374 = T384 ? T375 : 22'h0;
  assign T375 = T376;
  assign T376 = {R382, R377};
  assign T378 = T379 ? meta_io_resp_3_coh_state : R377;
  assign T379 = s1_clk_en & T380;
  assign T380 = s1_replaced_way_en[2'h3:2'h3];
  assign s1_replaced_way_en = 1'h1 << T381;
  assign T381 = R358[1'h1:1'h0];
  assign T383 = T379 ? meta_io_resp_3_tag : R382;
  assign T384 = s2_replaced_way_en[2'h3:2'h3];
  assign T385 = T396 | T386;
  assign T386 = T395 ? T387 : 22'h0;
  assign T387 = T388;
  assign T388 = {R393, R389};
  assign T390 = T391 ? meta_io_resp_2_coh_state : R389;
  assign T391 = s1_clk_en & T392;
  assign T392 = s1_replaced_way_en[2'h2:2'h2];
  assign T394 = T391 ? meta_io_resp_2_tag : R393;
  assign T395 = s2_replaced_way_en[2'h2:2'h2];
  assign T396 = T407 | T397;
  assign T397 = T406 ? T398 : 22'h0;
  assign T398 = T399;
  assign T399 = {R404, R400};
  assign T401 = T402 ? meta_io_resp_1_coh_state : R400;
  assign T402 = s1_clk_en & T403;
  assign T403 = s1_replaced_way_en[1'h1:1'h1];
  assign T405 = T402 ? meta_io_resp_1_tag : R404;
  assign T406 = s2_replaced_way_en[1'h1:1'h1];
  assign T407 = T416 ? T408 : 22'h0;
  assign T408 = T409;
  assign T409 = {R414, R410};
  assign T411 = T412 ? meta_io_resp_0_coh_state : R410;
  assign T412 = s1_clk_en & T413;
  assign T413 = s1_replaced_way_en[1'h0:1'h0];
  assign T415 = T412 ? meta_io_resp_0_tag : R414;
  assign T416 = s2_replaced_way_en[1'h0:1'h0];
  assign T417 = T44;
  assign T418 = s2_tag_match ? T420 : T419;
  assign T419 = T373[5'h15:2'h2];
  assign T420 = T419;
  assign T421 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T422 = s2_recycle ? s2_req_kill : T423;
  assign T423 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T424;
  assign T424 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T425 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T426 = s2_recycle ? s2_req_tag : T427;
  assign T427 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T428;
  assign T428 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T429 = s2_nack_hit ? 1'h0 : T430;
  assign T430 = T452 & T431;
  assign T431 = T439 | T432;
  assign T432 = T436 | T433;
  assign T433 = T435 | T434;
  assign T434 = s2_req_cmd == 5'h4;
  assign T435 = s2_req_cmd[2'h3:2'h3];
  assign T436 = T438 | T437;
  assign T437 = s2_req_cmd == 5'h7;
  assign T438 = s2_req_cmd == 5'h1;
  assign T439 = T449 | T440;
  assign T440 = T444 | T441;
  assign T441 = T443 | T442;
  assign T442 = s2_req_cmd == 5'h4;
  assign T443 = s2_req_cmd[2'h3:2'h3];
  assign T444 = T446 | T445;
  assign T445 = s2_req_cmd == 5'h7;
  assign T446 = T448 | T447;
  assign T447 = s2_req_cmd == 5'h6;
  assign T448 = s2_req_cmd == 5'h0;
  assign T449 = T451 | T450;
  assign T450 = s2_req_cmd == 5'h3;
  assign T451 = s2_req_cmd == 5'h2;
  assign T452 = s2_valid_masked & T453;
  assign T453 = s2_hit ^ 1'h1;
  assign T454 = io_mem_probe_valid & T455;
  assign T455 = lrsc_valid ^ 1'h1;
  assign io_mem_release_bits_data = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_voluntary = releaseArb_io_out_bits_voluntary;
  assign io_mem_release_bits_r_type = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_client_xact_id = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_addr_block = releaseArb_io_out_bits_addr_block;
  assign io_mem_release_bits_addr_beat = releaseArb_io_out_bits_addr_beat;
  assign io_mem_release_valid = releaseArb_io_out_valid;
  assign io_mem_probe_ready = T456;
  assign T456 = prober_io_req_ready & T457;
  assign T457 = lrsc_valid ^ 1'h1;
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_data = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_union = mshrs_io_mem_req_bits_union;
  assign io_mem_acquire_bits_a_type = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_is_builtin_type = mshrs_io_mem_req_bits_is_builtin_type;
  assign io_mem_acquire_bits_addr_beat = mshrs_io_mem_req_bits_addr_beat;
  assign io_mem_acquire_bits_client_xact_id = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_block = mshrs_io_mem_req_bits_addr_block;
  assign io_mem_acquire_valid = mshrs_io_mem_req_valid;
  assign io_ptw_req_bits_fetch = dtlb_io_ptw_req_bits_fetch;
  assign io_ptw_req_bits_store = dtlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_prv = dtlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_addr = dtlb_io_ptw_req_bits_addr;
  assign io_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_ordered = T458;
  assign T458 = T460 & T459;
  assign T459 = s2_valid ^ 1'h1;
  assign T460 = mshrs_io_fence_rdy & T461;
  assign T461 = s1_valid ^ 1'h1;
  assign io_cpu_xcpt_pf_st = T462;
  assign T462 = s1_write & dtlb_io_resp_xcpt_st;
  assign io_cpu_xcpt_pf_ld = T463;
  assign T463 = s1_read & dtlb_io_resp_xcpt_ld;
  assign io_cpu_xcpt_ma_st = T464;
  assign T464 = s1_write & misaligned;
  assign misaligned = T469 | T465;
  assign T465 = T468 & T466;
  assign T466 = T467 != 3'h0;
  assign T467 = s1_req_addr[2'h2:1'h0];
  assign T468 = s1_req_typ == 3'h3;
  assign T469 = T476 | T470;
  assign T470 = T473 & T471;
  assign T471 = T472 != 2'h0;
  assign T472 = s1_req_addr[1'h1:1'h0];
  assign T473 = T475 | T474;
  assign T474 = s1_req_typ == 3'h6;
  assign T475 = s1_req_typ == 3'h2;
  assign T476 = T479 & T477;
  assign T477 = T478 != 1'h0;
  assign T478 = s1_req_addr[1'h0:1'h0];
  assign T479 = T481 | T480;
  assign T480 = s1_req_typ == 3'h5;
  assign T481 = s1_req_typ == 3'h1;
  assign io_cpu_xcpt_ma_ld = T482;
  assign T482 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T483;
  assign T483 = s1_replay & s1_read;
  assign io_cpu_resp_bits_store_data = T484;
  assign T484 = cache_pass ? cache_resp_bits_store_data : uncache_resp_bits_store_data;
  assign uncache_resp_bits_store_data = mshrs_io_resp_bits_store_data;
  assign cache_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_data_word_bypass = T485;
  assign T485 = {T490, T486};
  assign T486 = T489 ? T488 : T487;
  assign T487 = s2_data_word[5'h1f:1'h0];
  assign T488 = s2_data_word[6'h3f:6'h20];
  assign T489 = s2_req_addr[2'h2:2'h2];
  assign T490 = T502 ? T492 : T491;
  assign T491 = s2_data_word[6'h3f:6'h20];
  assign T492 = 32'h0 - T604;
  assign T604 = {31'h0, T493};
  assign T493 = T495 & T494;
  assign T494 = T486[5'h1f:5'h1f];
  assign T495 = T497 | T496;
  assign T496 = s2_req_typ == 3'h3;
  assign T497 = T499 | T498;
  assign T498 = s2_req_typ == 3'h2;
  assign T499 = T501 | T500;
  assign T500 = s2_req_typ == 3'h1;
  assign T501 = s2_req_typ == 3'h0;
  assign T502 = T504 | T503;
  assign T503 = s2_req_typ == 3'h6;
  assign T504 = s2_req_typ == 3'h2;
  assign io_cpu_resp_bits_has_data = T505;
  assign T505 = cache_pass ? cache_resp_bits_has_data : uncache_resp_bits_has_data;
  assign uncache_resp_bits_has_data = mshrs_io_resp_bits_has_data;
  assign cache_resp_bits_has_data = T506;
  assign T506 = T510 | T507;
  assign T507 = T509 | T508;
  assign T508 = s2_req_cmd == 5'h4;
  assign T509 = s2_req_cmd[2'h3:2'h3];
  assign T510 = T512 | T511;
  assign T511 = s2_req_cmd == 5'h7;
  assign T512 = T514 | T513;
  assign T513 = s2_req_cmd == 5'h6;
  assign T514 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_replay = T515;
  assign T515 = cache_pass ? cache_resp_bits_replay : uncache_resp_bits_replay;
  assign uncache_resp_bits_replay = mshrs_io_resp_bits_replay;
  assign cache_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T516;
  assign T516 = cache_pass ? cache_resp_bits_nack : uncache_resp_bits_nack;
  assign uncache_resp_bits_nack = mshrs_io_resp_bits_nack;
  assign cache_resp_bits_nack = T517;
  assign T517 = s2_valid & s2_nack;
  assign io_cpu_resp_bits_data = T518;
  assign T518 = cache_pass ? cache_resp_bits_data : uncache_resp_bits_data;
  assign uncache_resp_bits_data = mshrs_io_resp_bits_data;
  assign cache_resp_bits_data = T519;
  assign T519 = T520 | T605;
  assign T605 = {63'h0, s2_sc_fail};
  assign T520 = {T539, T521};
  assign T521 = s2_sc ? 8'h0 : T522;
  assign T522 = T538 ? T537 : T523;
  assign T523 = T524[3'h7:1'h0];
  assign T524 = {T529, T525};
  assign T525 = T528 ? T527 : T526;
  assign T526 = T485[4'hf:1'h0];
  assign T527 = T485[5'h1f:5'h10];
  assign T528 = s2_req_addr[1'h1:1'h1];
  assign T529 = T534 ? T531 : T530;
  assign T530 = T485[6'h3f:5'h10];
  assign T531 = 48'h0 - T606;
  assign T606 = {47'h0, T532};
  assign T532 = T495 & T533;
  assign T533 = T525[4'hf:4'hf];
  assign T534 = T536 | T535;
  assign T535 = s2_req_typ == 3'h5;
  assign T536 = s2_req_typ == 3'h1;
  assign T537 = T524[4'hf:4'h8];
  assign T538 = s2_req_addr[1'h0:1'h0];
  assign T539 = T544 ? T541 : T540;
  assign T540 = T524[6'h3f:4'h8];
  assign T541 = 56'h0 - T607;
  assign T607 = {55'h0, T542};
  assign T542 = T495 & T543;
  assign T543 = T521[3'h7:3'h7];
  assign T544 = s2_sc | T545;
  assign T545 = T547 | T546;
  assign T546 = s2_req_typ == 3'h4;
  assign T547 = s2_req_typ == 3'h0;
  assign io_cpu_resp_bits_typ = T548;
  assign T548 = cache_pass ? cache_resp_bits_typ : uncache_resp_bits_typ;
  assign uncache_resp_bits_typ = mshrs_io_resp_bits_typ;
  assign cache_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_cmd = T549;
  assign T549 = cache_pass ? cache_resp_bits_cmd : uncache_resp_bits_cmd;
  assign uncache_resp_bits_cmd = mshrs_io_resp_bits_cmd;
  assign cache_resp_bits_cmd = s2_req_cmd;
  assign io_cpu_resp_bits_tag = T550;
  assign T550 = cache_pass ? cache_resp_bits_tag : uncache_resp_bits_tag;
  assign uncache_resp_bits_tag = mshrs_io_resp_bits_tag;
  assign cache_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_addr = T551;
  assign T551 = cache_pass ? cache_resp_bits_addr : uncache_resp_bits_addr;
  assign uncache_resp_bits_addr = mshrs_io_resp_bits_addr;
  assign cache_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_valid = T552;
  assign T552 = cache_pass ? cache_resp_valid : uncache_resp_valid;
  assign uncache_resp_valid = mshrs_io_resp_valid;
  assign cache_resp_valid = T553;
  assign T553 = T555 & T554;
  assign T554 = s2_data_correctable ^ 1'h1;
  assign T555 = s2_replay | T556;
  assign T556 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T557;
  assign T557 = block_miss ? 1'h0 : T558;
  assign T558 = T565 ? 1'h0 : T559;
  assign T559 = T564 ? 1'h0 : T560;
  assign T560 = T561 == 1'h0;
  assign T561 = T563 & T562;
  assign T562 = io_cpu_req_bits_phys ^ 1'h1;
  assign T563 = dtlb_io_req_ready ^ 1'h1;
  assign T564 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T565 = readArb_io_in_3_ready ^ 1'h1;
  assign T608 = reset ? 1'h0 : T566;
  assign T566 = T567 & s2_nack_miss;
  assign T567 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_addr_beat( wbArb_io_out_bits_addr_beat ),
       .io_req_bits_addr_block( wbArb_io_out_bits_addr_block ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_req_bits_voluntary( wbArb_io_out_bits_voluntary ),
       .io_req_bits_data( wbArb_io_out_bits_data ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( s2_data_corrected ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr_beat( wb_io_release_bits_addr_beat ),
       .io_release_bits_addr_block( wb_io_release_bits_addr_block ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_r_type( wb_io_release_bits_r_type ),
       .io_release_bits_voluntary( wb_io_release_bits_voluntary ),
       .io_release_bits_data( wb_io_release_bits_data )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T454 ),
       .io_req_bits_addr_block( io_mem_probe_bits_addr_block ),
       .io_req_bits_p_type( io_mem_probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr_beat( prober_io_rep_bits_addr_beat ),
       .io_rep_bits_addr_block( prober_io_rep_bits_addr_block ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_rep_bits_voluntary( prober_io_rep_bits_voluntary ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( prober_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( prober_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_wb_req_bits_voluntary( prober_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_data( prober_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_block_state_state( T44 )
  );
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T429 ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_data( s2_req_data ),
       .io_req_bits_tag_match( s2_tag_match ),
       .io_req_bits_old_meta_tag( T418 ),
       .io_req_bits_old_meta_coh_state( T371 ),
       .io_req_bits_way_en( T354 ),
       .io_resp_ready( T353 ),
       .io_resp_valid( mshrs_io_resp_valid ),
       .io_resp_bits_addr( mshrs_io_resp_bits_addr ),
       .io_resp_bits_tag( mshrs_io_resp_bits_tag ),
       .io_resp_bits_cmd( mshrs_io_resp_bits_cmd ),
       .io_resp_bits_typ( mshrs_io_resp_bits_typ ),
       .io_resp_bits_data( mshrs_io_resp_bits_data ),
       .io_resp_bits_nack( mshrs_io_resp_bits_nack ),
       .io_resp_bits_replay( mshrs_io_resp_bits_replay ),
       .io_resp_bits_has_data( mshrs_io_resp_bits_has_data ),
       //.io_resp_bits_data_word_bypass(  )
       .io_resp_bits_store_data( mshrs_io_resp_bits_store_data ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( io_mem_acquire_ready ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( mshrs_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( mshrs_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_is_builtin_type( mshrs_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( mshrs_io_mem_req_bits_union ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_refill_way_en( mshrs_io_refill_way_en ),
       .io_refill_addr( mshrs_io_refill_addr ),
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_mem_grant_valid( T352 ),
       .io_mem_grant_bits_addr_beat( FlowThroughSerializer_io_out_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( FlowThroughSerializer_io_out_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( FlowThroughSerializer_io_out_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( FlowThroughSerializer_io_out_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( FlowThroughSerializer_io_out_bits_g_type ),
       .io_mem_grant_bits_data( FlowThroughSerializer_io_out_bits_data ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( mshrs_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( mshrs_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_wb_req_bits_voluntary( mshrs_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_data( mshrs_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T337 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T336 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_req_bits_store( s1_write ),
       .io_resp_miss( dtlb_io_resp_miss ),
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       //.io_resp_hit_idx(  )
       .io_ptw_req_ready( io_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( dtlb_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( dtlb_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( dtlb_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( dtlb_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( io_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_ptw_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( io_ptw_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( io_ptw_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( io_ptw_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( io_ptw_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( io_ptw_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( io_ptw_resp_bits_pte_v ),
       .io_ptw_status_sd( io_ptw_status_sd ),
       .io_ptw_status_zero2( io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( io_ptw_status_zero1 ),
       .io_ptw_status_vm( io_ptw_status_vm ),
       .io_ptw_status_mprv( io_ptw_status_mprv ),
       .io_ptw_status_xs( io_ptw_status_xs ),
       .io_ptw_status_fs( io_ptw_status_fs ),
       .io_ptw_status_prv3( io_ptw_status_prv3 ),
       .io_ptw_status_ie3( io_ptw_status_ie3 ),
       .io_ptw_status_prv2( io_ptw_status_prv2 ),
       .io_ptw_status_ie2( io_ptw_status_ie2 ),
       .io_ptw_status_prv1( io_ptw_status_prv1 ),
       .io_ptw_status_ie1( io_ptw_status_ie1 ),
       .io_ptw_status_prv( io_ptw_status_prv ),
       .io_ptw_status_ie( io_ptw_status_ie ),
       .io_ptw_invalidate( io_ptw_invalidate )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_3_tag( meta_io_resp_3_tag ),
       .io_resp_3_coh_state( meta_io_resp_3_coh_state ),
       .io_resp_2_tag( meta_io_resp_2_tag ),
       .io_resp_2_coh_state( meta_io_resp_2_coh_state ),
       .io_resp_1_tag( meta_io_resp_1_tag ),
       .io_resp_1_coh_state( meta_io_resp_1_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state )
  );
  Arbiter_0 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T602 ),
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T601 ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx )
       //.io_chosen(  )
  );
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T326 ),
       .io_resp_3( data_io_resp_3 ),
       .io_resp_2( data_io_resp_2 ),
       .io_resp_1( data_io_resp_1 ),
       .io_resp_0( data_io_resp_0 )
  );
  Arbiter_2 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 4'hf ),
       .io_in_3_bits_addr( T600 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 4'hf ),
       .io_in_1_bits_addr( T599 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 4'hf ),
       .io_in_0_bits_addr( T598 ),
       .io_out_ready( T324 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_3 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T314 ),
       .io_in_1_bits_way_en( mshrs_io_refill_way_en ),
       .io_in_1_bits_addr( mshrs_io_refill_addr ),
       .io_in_1_bits_wmask( 2'h3 ),
       .io_in_1_bits_data( FlowThroughSerializer_io_out_bits_data ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T597 ),
       .io_in_0_bits_wmask( rowWMask ),
       .io_in_0_bits_data( T311 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T596 ),
       .io_cmd( s2_req_cmd ),
       .io_typ( s2_req_typ ),
       .io_lhs( T577 ),
       .io_rhs( s2_req_data ),
       .io_out( amoalu_io_out )
  );
  LockingArbiter_0 releaseArb(.clk(clk), .reset(reset),
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr_beat( prober_io_rep_bits_addr_beat ),
       .io_in_1_bits_addr_block( prober_io_rep_bits_addr_block ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_1_bits_voluntary( prober_io_rep_bits_voluntary ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr_beat( wb_io_release_bits_addr_beat ),
       .io_in_0_bits_addr_block( wb_io_release_bits_addr_block ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_in_0_bits_voluntary( wb_io_release_bits_voluntary ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_out_ready( io_mem_release_ready ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr_beat( releaseArb_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( releaseArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type ),
       .io_out_bits_voluntary( releaseArb_io_out_bits_voluntary ),
       .io_out_bits_data( releaseArb_io_out_bits_data )
       //.io_chosen(  )
  );
  FlowThroughSerializer FlowThroughSerializer(
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_in_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_in_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_in_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_in_bits_g_type( io_mem_grant_bits_g_type ),
       .io_in_bits_data( io_mem_grant_bits_data ),
       .io_out_ready( T8 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       .io_out_bits_addr_beat( FlowThroughSerializer_io_out_bits_addr_beat ),
       .io_out_bits_client_xact_id( FlowThroughSerializer_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( FlowThroughSerializer_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( FlowThroughSerializer_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( FlowThroughSerializer_io_out_bits_g_type ),
       .io_out_bits_data( FlowThroughSerializer_io_out_bits_data )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_4 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_addr_beat( mshrs_io_wb_req_bits_addr_beat ),
       .io_in_1_bits_addr_block( mshrs_io_wb_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_1_bits_voluntary( mshrs_io_wb_req_bits_voluntary ),
       .io_in_1_bits_data( mshrs_io_wb_req_bits_data ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_addr_beat( prober_io_wb_req_bits_addr_beat ),
       .io_in_0_bits_addr_block( prober_io_wb_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_in_0_bits_voluntary( prober_io_wb_req_bits_voluntary ),
       .io_in_0_bits_data( prober_io_wb_req_bits_data ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_addr_beat( wbArb_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( wbArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_out_bits_voluntary( wbArb_io_out_bits_voluntary ),
       .io_out_bits_data( wbArb_io_out_bits_data ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "DCache exception occurred - cache response not killed.");
    $finish;
  end
// synthesis translate_on
`endif
    R4 <= T5;
    if(T138) begin
      s2_req_data <= s1_req_data;
    end else if(T21) begin
      s2_req_data <= T19;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T20;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T30) begin
      s2_recycle_next <= s2_recycle_ecc;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T31;
    end
    if(s1_clk_en) begin
      R48 <= meta_io_resp_3_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T572;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T571;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T573;
    end
    if(s1_clk_en) begin
      R92 <= meta_io_resp_2_coh_state;
    end
    if(s1_clk_en) begin
      R98 <= meta_io_resp_1_coh_state;
    end
    if(s1_clk_en) begin
      R103 <= meta_io_resp_0_coh_state;
    end
    if(reset) begin
      R129 <= 1'h0;
    end else begin
      R129 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(reset) begin
      s1_recycled <= 1'h0;
    end else if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R145 <= T578;
    if(T153) begin
      R150 <= T152;
    end
    R162 <= T580;
    if(T170) begin
      R167 <= T169;
    end
    R176 <= T582;
    if(T184) begin
      R181 <= T183;
    end
    R189 <= T584;
    if(T197) begin
      R194 <= T196;
    end
    if(T288) begin
      s2_store_bypass_data <= T201;
    end
    if(T204) begin
      s4_req_data <= s3_req_data;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T205;
    end
    if(T220) begin
      lrsc_addr <= T219;
    end
    if(T234) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_invalidate_lr) begin
      lrsc_count <= 5'h0;
    end else if(T242) begin
      lrsc_count <= 5'h0;
    end else if(T240) begin
      lrsc_count <= 5'h1f;
    end else if(lrsc_valid) begin
      lrsc_count <= T239;
    end
    s3_req_data <= T589;
    if(T249) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T249) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T204) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T204) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T288) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T249) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    if(s1_clk_en) begin
      R355 <= T357;
    end
    if(reset) begin
      R358 <= 16'h1;
    end else if(T369) begin
      R358 <= T360;
    end
    if(T379) begin
      R377 <= meta_io_resp_3_coh_state;
    end
    if(T379) begin
      R382 <= meta_io_resp_3_tag;
    end
    if(T391) begin
      R389 <= meta_io_resp_2_coh_state;
    end
    if(T391) begin
      R393 <= meta_io_resp_2_tag;
    end
    if(T402) begin
      R400 <= meta_io_resp_1_coh_state;
    end
    if(T402) begin
      R404 <= meta_io_resp_1_tag;
    end
    if(T412) begin
      R410 <= meta_io_resp_0_coh_state;
    end
    if(T412) begin
      R414 <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T566;
    end
  end
endmodule

module RRArbiter_2(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [26:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_prv,
    input  io_in_1_bits_store,
    input  io_in_1_bits_fetch,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [26:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_prv,
    input  io_in_0_bits_store,
    input  io_in_0_bits_fetch,
    input  io_out_ready,
    output io_out_valid,
    output[26:0] io_out_bits_addr,
    output[1:0] io_out_bits_prv,
    output io_out_bits_store,
    output io_out_bits_fetch,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T28;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[1:0] T8;
  wire[26:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T28 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_fetch = T5;
  assign T5 = T6 ? io_in_1_bits_fetch : io_in_0_bits_fetch;
  assign T6 = chosen;
  assign io_out_bits_store = T7;
  assign T7 = T6 ? io_in_1_bits_store : io_in_0_bits_store;
  assign io_out_bits_prv = T8;
  assign T8 = T6 ? io_in_1_bits_prv : io_in_0_bits_prv;
  assign io_out_bits_addr = T9;
  assign T9 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T10;
  assign T10 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = T19 | T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = T17 | T15;
  assign T15 = io_in_1_valid & T16;
  assign T16 = last_grant < 1'h1;
  assign T17 = io_in_0_valid & T18;
  assign T18 = last_grant < 1'h0;
  assign T19 = last_grant < 1'h0;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = T25 | T22;
  assign T22 = T23 ^ 1'h1;
  assign T23 = T24 | io_in_0_valid;
  assign T24 = T17 | T15;
  assign T25 = T27 & T26;
  assign T26 = last_grant < 1'h1;
  assign T27 = T17 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [26:0] io_requestor_1_req_bits_addr,
    input [1:0] io_requestor_1_req_bits_prv,
    input  io_requestor_1_req_bits_store,
    input  io_requestor_1_req_bits_fetch,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[19:0] io_requestor_1_resp_bits_pte_ppn,
    output[2:0] io_requestor_1_resp_bits_pte_reserved_for_software,
    output io_requestor_1_resp_bits_pte_d,
    output io_requestor_1_resp_bits_pte_r,
    output[3:0] io_requestor_1_resp_bits_pte_typ,
    output io_requestor_1_resp_bits_pte_v,
    output io_requestor_1_status_sd,
    output[30:0] io_requestor_1_status_zero2,
    output io_requestor_1_status_sd_rv32,
    output[8:0] io_requestor_1_status_zero1,
    output[4:0] io_requestor_1_status_vm,
    output io_requestor_1_status_mprv,
    output[1:0] io_requestor_1_status_xs,
    output[1:0] io_requestor_1_status_fs,
    output[1:0] io_requestor_1_status_prv3,
    output io_requestor_1_status_ie3,
    output[1:0] io_requestor_1_status_prv2,
    output io_requestor_1_status_ie2,
    output[1:0] io_requestor_1_status_prv1,
    output io_requestor_1_status_ie1,
    output[1:0] io_requestor_1_status_prv,
    output io_requestor_1_status_ie,
    output io_requestor_1_invalidate,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [26:0] io_requestor_0_req_bits_addr,
    input [1:0] io_requestor_0_req_bits_prv,
    input  io_requestor_0_req_bits_store,
    input  io_requestor_0_req_bits_fetch,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[19:0] io_requestor_0_resp_bits_pte_ppn,
    output[2:0] io_requestor_0_resp_bits_pte_reserved_for_software,
    output io_requestor_0_resp_bits_pte_d,
    output io_requestor_0_resp_bits_pte_r,
    output[3:0] io_requestor_0_resp_bits_pte_typ,
    output io_requestor_0_resp_bits_pte_v,
    output io_requestor_0_status_sd,
    output[30:0] io_requestor_0_status_zero2,
    output io_requestor_0_status_sd_rv32,
    output[8:0] io_requestor_0_status_zero1,
    output[4:0] io_requestor_0_status_vm,
    output io_requestor_0_status_mprv,
    output[1:0] io_requestor_0_status_xs,
    output[1:0] io_requestor_0_status_fs,
    output[1:0] io_requestor_0_status_prv3,
    output io_requestor_0_status_ie3,
    output[1:0] io_requestor_0_status_prv2,
    output io_requestor_0_status_ie2,
    output[1:0] io_requestor_0_status_prv1,
    output io_requestor_0_status_ie1,
    output[1:0] io_requestor_0_status_prv,
    output io_requestor_0_status_ie,
    output io_requestor_0_invalidate,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[39:0] io_mem_req_bits_addr,
    //output[8:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_kill,
    output io_mem_req_bits_phys,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [39:0] io_mem_resp_bits_addr,
    input [8:0] io_mem_resp_bits_tag,
    input [4:0] io_mem_resp_bits_cmd,
    input [2:0] io_mem_resp_bits_typ,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_word_bypass,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [8:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_invalidate_lr
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_status_sd,
    input [30:0] io_dpath_status_zero2,
    input  io_dpath_status_sd_rv32,
    input [8:0] io_dpath_status_zero1,
    input [4:0] io_dpath_status_vm,
    input  io_dpath_status_mprv,
    input [1:0] io_dpath_status_xs,
    input [1:0] io_dpath_status_fs,
    input [1:0] io_dpath_status_prv3,
    input  io_dpath_status_ie3,
    input [1:0] io_dpath_status_prv2,
    input  io_dpath_status_ie2,
    input [1:0] io_dpath_status_prv1,
    input  io_dpath_status_ie1,
    input [1:0] io_dpath_status_prv,
    input  io_dpath_status_ie
);

  wire T0;
  reg [2:0] state;
  wire[2:0] T232;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [1:0] count;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire pte_cache_hit;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[1:0] T26;
  reg  R27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T233;
  wire[1:0] T234;
  wire T235;
  wire[2:0] T36;
  wire T236;
  wire[1:0] T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire T44;
  reg [2:0] R45;
  wire[2:0] T46;
  wire[2:0] T47;
  wire[2:0] T48;
  wire[2:0] T49;
  wire[5:0] T50;
  wire[1:0] T51;
  wire T52;
  wire[1:0] T237;
  wire T238;
  wire[1:0] T239;
  wire[1:0] T240;
  wire T241;
  wire T242;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire[2:0] T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[3:0] T70;
  wire T71;
  wire T72;
  reg  R73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg  R78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire T86;
  wire[31:0] pte_addr;
  wire[28:0] T87;
  wire[28:0] T88;
  wire[8:0] vpn_idx;
  wire[8:0] T89;
  wire[8:0] T90;
  wire[8:0] T91;
  reg [26:0] r_req_addr;
  wire[26:0] T92;
  wire T93;
  wire[8:0] T94;
  wire[17:0] T95;
  wire T96;
  wire[1:0] T97;
  wire[8:0] T98;
  wire[26:0] T99;
  wire T100;
  reg [19:0] r_pte_ppn;
  wire[19:0] T101;
  wire[19:0] T102;
  wire[19:0] T103;
  wire[19:0] T104;
  wire[19:0] T105;
  wire T106;
  wire T107;
  wire set_dirty_bit;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg  r_req_store;
  wire T112;
  wire T113;
  wire T114;
  wire perm_ok;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg  r_req_fetch;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  reg [1:0] r_req_prv;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire[19:0] pte_cache_data;
  wire[19:0] T150;
  wire[19:0] T151;
  reg [19:0] T152 [2:0];
  wire[19:0] T153;
  wire T154;
  wire T155;
  wire[1:0] T156;
  wire T157;
  wire[19:0] T158;
  wire[19:0] T159;
  wire[19:0] T160;
  wire T161;
  wire[19:0] T162;
  wire[19:0] T163;
  wire T164;
  wire[31:0] T165;
  reg [31:0] T166 [2:0];
  wire[31:0] T167;
  wire T168;
  wire T169;
  wire[1:0] T170;
  wire T171;
  wire[31:0] T172;
  wire T173;
  wire[31:0] T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[2:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire[63:0] T243;
  wire[29:0] T198;
  wire[29:0] T199;
  wire[5:0] T200;
  wire[4:0] T201;
  wire pte_wdata_v;
  wire[3:0] pte_wdata_typ;
  wire pte_wdata_r;
  wire[23:0] T202;
  wire[3:0] T203;
  wire pte_wdata_d;
  wire[2:0] pte_wdata_reserved_for_software;
  wire[19:0] pte_wdata_ppn;
  wire[4:0] T204;
  wire T205;
  wire[39:0] T244;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  reg  r_pte_v;
  wire T210;
  reg [3:0] r_pte_typ;
  wire[3:0] T211;
  reg  r_pte_r;
  wire T212;
  reg  r_pte_d;
  wire T213;
  reg [2:0] r_pte_reserved_for_software;
  wire[2:0] T214;
  wire[2:0] T215;
  wire[19:0] T245;
  wire[27:0] resp_ppn;
  wire[27:0] T216;
  wire[27:0] T217;
  wire[17:0] T218;
  wire[9:0] T219;
  wire[27:0] T220;
  wire[8:0] T221;
  wire[18:0] T222;
  wire T223;
  wire[1:0] T224;
  wire[27:0] r_resp_ppn;
  wire T225;
  wire resp_err;
  wire T226;
  wire T227;
  reg  r_req_dest;
  wire T228;
  wire resp_val;
  wire T229;
  wire[19:0] T246;
  wire T230;
  wire T231;
  wire arb_io_in_1_ready;
  wire arb_io_in_0_ready;
  wire arb_io_out_valid;
  wire[26:0] arb_io_out_bits_addr;
  wire[1:0] arb_io_out_bits_prv;
  wire arb_io_out_bits_store;
  wire arb_io_out_bits_fetch;
  wire arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    R27 = {1{$random}};
    R45 = {1{$random}};
    R73 = {1{$random}};
    R78 = {1{$random}};
    r_req_addr = {1{$random}};
    r_pte_ppn = {1{$random}};
    r_req_store = {1{$random}};
    r_req_fetch = {1{$random}};
    r_req_prv = {1{$random}};
    for (initvar = 0; initvar < 3; initvar = initvar+1)
      T152[initvar] = {1{$random}};
    for (initvar = 0; initvar < 3; initvar = initvar+1)
      T166[initvar] = {1{$random}};
    r_pte_v = {1{$random}};
    r_pte_typ = {1{$random}};
    r_pte_r = {1{$random}};
    r_pte_d = {1{$random}};
    r_pte_reserved_for_software = {1{$random}};
    r_req_dest = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_invalidate_lr = {1{$random}};
//  assign io_mem_req_bits_tag = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = state == 3'h0;
  assign T232 = reset ? 3'h0 : T1;
  assign T1 = T197 ? 3'h0 : T2;
  assign T2 = T196 ? 3'h0 : T3;
  assign T3 = T195 ? 3'h1 : T4;
  assign T4 = T193 ? 3'h3 : T5;
  assign T5 = T191 ? 3'h4 : T6;
  assign T6 = T188 ? T187 : T7;
  assign T7 = T182 ? 3'h1 : T8;
  assign T8 = T181 ? 3'h6 : T9;
  assign T9 = T179 ? 3'h1 : T10;
  assign T10 = T176 ? 3'h2 : T11;
  assign T11 = T15 ? 3'h1 : T12;
  assign T12 = T13 ? 3'h1 : state;
  assign T13 = T14 & arb_io_out_valid;
  assign T14 = 3'h0 == state;
  assign T15 = T175 & T16;
  assign T16 = pte_cache_hit & T17;
  assign T17 = count < 2'h2;
  assign T18 = T182 ? T22 : T19;
  assign T19 = T15 ? T21 : T20;
  assign T20 = T14 ? 2'h0 : count;
  assign T21 = count + 2'h1;
  assign T22 = count + 2'h1;
  assign pte_cache_hit = T23 != 3'h0;
  assign T23 = T83 & T24;
  assign T24 = T25;
  assign T25 = {R78, T26};
  assign T26 = {R73, R27};
  assign T28 = T72 ? 1'h0 : T29;
  assign T29 = T30 ? 1'h1 : R27;
  assign T30 = T65 & T31;
  assign T31 = T32[1'h0:1'h0];
  assign T32 = 1'h1 << T33;
  assign T33 = T34;
  assign T34 = T64 ? T37 : T233;
  assign T233 = T236 ? 1'h0 : T234;
  assign T234 = T235 ? 1'h1 : 2'h2;
  assign T235 = T36[1'h1:1'h1];
  assign T36 = ~ T24;
  assign T236 = T36[1'h0:1'h0];
  assign T37 = T38[1'h1:1'h0];
  assign T38 = {T62, T39};
  assign T39 = T44 & T40;
  assign T40 = T41 - 1'h1;
  assign T41 = 1'h1 << T42;
  assign T42 = T43 + 2'h1;
  assign T43 = T62 - T62;
  assign T44 = R45 >> T62;
  assign T46 = T60 ? T47 : R45;
  assign T47 = T55 | T48;
  assign T48 = T54 ? 3'h0 : T49;
  assign T49 = T50[2'h2:1'h0];
  assign T50 = 3'h1 << T51;
  assign T51 = {1'h1, T52};
  assign T52 = T237[1'h1:1'h1];
  assign T237 = {T242, T238};
  assign T238 = T239[1'h1:1'h1];
  assign T239 = T241 | T240;
  assign T240 = T23[1'h1:1'h0];
  assign T241 = T23[2'h2:2'h2];
  assign T242 = T241 != 1'h0;
  assign T54 = T237[1'h0:1'h0];
  assign T55 = T57 & T56;
  assign T56 = ~ T49;
  assign T57 = T59 | T58;
  assign T58 = T52 ? 3'h0 : 3'h2;
  assign T59 = R45 & 3'h5;
  assign T60 = pte_cache_hit & T61;
  assign T61 = state == 3'h1;
  assign T62 = {1'h1, T63};
  assign T63 = R45[1'h1:1'h1];
  assign T64 = T24 == 3'h7;
  assign T65 = T67 & T66;
  assign T66 = pte_cache_hit ^ 1'h1;
  assign T67 = io_mem_resp_valid & T68;
  assign T68 = T71 & T69;
  assign T69 = T70 < 4'h2;
  assign T70 = io_mem_resp_bits_data[3'h4:1'h1];
  assign T71 = io_mem_resp_bits_data[1'h0:1'h0];
  assign T72 = reset | io_dpath_invalidate;
  assign T74 = T72 ? 1'h0 : T75;
  assign T75 = T76 ? 1'h1 : R73;
  assign T76 = T65 & T77;
  assign T77 = T32[1'h1:1'h1];
  assign T79 = T72 ? 1'h0 : T80;
  assign T80 = T81 ? 1'h1 : R78;
  assign T81 = T65 & T82;
  assign T82 = T32[2'h2:2'h2];
  assign T83 = T84;
  assign T84 = {T173, T85};
  assign T85 = {T171, T86};
  assign T86 = T165 == pte_addr;
  assign pte_addr = T87 << 2'h3;
  assign T87 = T88;
  assign T88 = {r_pte_ppn, vpn_idx};
  assign vpn_idx = T100 ? T98 : T89;
  assign T89 = T96 ? T94 : T90;
  assign T90 = T91[4'h8:1'h0];
  assign T91 = r_req_addr >> 5'h12;
  assign T92 = T93 ? arb_io_out_bits_addr : r_req_addr;
  assign T93 = T0 & arb_io_out_valid;
  assign T94 = T95[4'h8:1'h0];
  assign T95 = r_req_addr >> 4'h9;
  assign T96 = T97[1'h0:1'h0];
  assign T97 = count;
  assign T98 = T99[4'h8:1'h0];
  assign T99 = r_req_addr >> 1'h0;
  assign T100 = T97[1'h1:1'h1];
  assign T101 = T15 ? pte_cache_data : T102;
  assign T102 = T106 ? T105 : T103;
  assign T103 = T93 ? T104 : r_pte_ppn;
  assign T104 = io_dpath_ptbr[5'h1f:4'hc];
  assign T105 = io_mem_resp_bits_data[5'h1d:4'ha];
  assign T106 = T148 & T107;
  assign T107 = set_dirty_bit ^ 1'h1;
  assign set_dirty_bit = perm_ok & T108;
  assign T108 = T113 | T109;
  assign T109 = r_req_store & T110;
  assign T110 = T111 ^ 1'h1;
  assign T111 = io_mem_resp_bits_data[3'h6:3'h6];
  assign T112 = T93 ? arb_io_out_bits_store : r_req_store;
  assign T113 = T114 ^ 1'h1;
  assign T114 = io_mem_resp_bits_data[3'h5:3'h5];
  assign perm_ok = T146 ? T134 : T115;
  assign T115 = r_req_fetch ? T127 : T116;
  assign T116 = r_req_store ? T121 : T117;
  assign T117 = T119 & T118;
  assign T118 = T70 < 4'h8;
  assign T119 = T71 & T120;
  assign T120 = 4'h2 <= T70;
  assign T121 = T123 & T122;
  assign T122 = T70[1'h0:1'h0];
  assign T123 = T125 & T124;
  assign T124 = T70 < 4'h8;
  assign T125 = T71 & T126;
  assign T126 = 4'h2 <= T70;
  assign T127 = T129 & T128;
  assign T128 = T70[1'h1:1'h1];
  assign T129 = T131 & T130;
  assign T130 = T70 < 4'h8;
  assign T131 = T71 & T132;
  assign T132 = 4'h2 <= T70;
  assign T133 = T93 ? arb_io_out_bits_fetch : r_req_fetch;
  assign T134 = r_req_fetch ? T142 : T135;
  assign T135 = r_req_store ? T138 : T136;
  assign T136 = T71 & T137;
  assign T137 = 4'h2 <= T70;
  assign T138 = T140 & T139;
  assign T139 = T70[1'h0:1'h0];
  assign T140 = T71 & T141;
  assign T141 = 4'h2 <= T70;
  assign T142 = T144 & T143;
  assign T143 = T70[1'h1:1'h1];
  assign T144 = T71 & T145;
  assign T145 = 4'h4 <= T70;
  assign T146 = r_req_prv[1'h0:1'h0];
  assign T147 = T93 ? arb_io_out_bits_prv : r_req_prv;
  assign T148 = io_mem_resp_valid & T149;
  assign T149 = state == 3'h2;
  assign pte_cache_data = T158 | T150;
  assign T150 = T157 ? T151 : 20'h0;
  assign T151 = T152[2'h2];
  assign T154 = T65 & T155;
  assign T155 = T156 < 2'h3;
  assign T156 = T34[1'h1:1'h0];
  assign T157 = T23[2'h2:2'h2];
  assign T158 = T162 | T159;
  assign T159 = T161 ? T160 : 20'h0;
  assign T160 = T152[2'h1];
  assign T161 = T23[1'h1:1'h1];
  assign T162 = T164 ? T163 : 20'h0;
  assign T163 = T152[2'h0];
  assign T164 = T23[1'h0:1'h0];
  assign T165 = T166[2'h0];
  assign T168 = T65 & T169;
  assign T169 = T170 < 2'h3;
  assign T170 = T34[1'h1:1'h0];
  assign T171 = T172 == pte_addr;
  assign T172 = T166[2'h1];
  assign T173 = T174 == pte_addr;
  assign T174 = T166[2'h2];
  assign T175 = 3'h1 == state;
  assign T176 = T175 & T177;
  assign T177 = T178 & io_mem_req_ready;
  assign T178 = T16 ^ 1'h1;
  assign T179 = T180 & io_mem_resp_bits_nack;
  assign T180 = 3'h2 == state;
  assign T181 = T180 & io_mem_resp_valid;
  assign T182 = T181 & T183;
  assign T183 = T185 & T184;
  assign T184 = count < 2'h2;
  assign T185 = T71 & T186;
  assign T186 = T70 < 4'h2;
  assign T187 = set_dirty_bit ? 3'h3 : 3'h5;
  assign T188 = T181 & T189;
  assign T189 = T71 & T190;
  assign T190 = 4'h2 <= T70;
  assign T191 = T192 & io_mem_req_ready;
  assign T192 = 3'h3 == state;
  assign T193 = T194 & io_mem_resp_bits_nack;
  assign T194 = 3'h4 == state;
  assign T195 = T194 & io_mem_resp_valid;
  assign T196 = 3'h5 == state;
  assign T197 = 3'h6 == state;
  assign io_mem_req_bits_data = T243;
  assign T243 = {34'h0, T198};
  assign T198 = T199;
  assign T199 = {T202, T200};
  assign T200 = {pte_wdata_r, T201};
  assign T201 = {pte_wdata_typ, pte_wdata_v};
  assign pte_wdata_v = 1'h0;
  assign pte_wdata_typ = 4'h0;
  assign pte_wdata_r = 1'h1;
  assign T202 = {pte_wdata_ppn, T203};
  assign T203 = {pte_wdata_reserved_for_software, pte_wdata_d};
  assign pte_wdata_d = r_req_store;
  assign pte_wdata_reserved_for_software = 3'h0;
  assign pte_wdata_ppn = 20'h0;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_cmd = T204;
  assign T204 = T205 ? 5'ha : 5'h0;
  assign T205 = state == 3'h3;
  assign io_mem_req_bits_addr = T244;
  assign T244 = {8'h0, pte_addr};
  assign io_mem_req_valid = T206;
  assign T206 = T15 ? 1'h0 : T207;
  assign T207 = T209 | T208;
  assign T208 = state == 3'h3;
  assign T209 = state == 3'h1;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_ie = io_dpath_status_ie;
  assign io_requestor_0_status_prv = io_dpath_status_prv;
  assign io_requestor_0_status_ie1 = io_dpath_status_ie1;
  assign io_requestor_0_status_prv1 = io_dpath_status_prv1;
  assign io_requestor_0_status_ie2 = io_dpath_status_ie2;
  assign io_requestor_0_status_prv2 = io_dpath_status_prv2;
  assign io_requestor_0_status_ie3 = io_dpath_status_ie3;
  assign io_requestor_0_status_prv3 = io_dpath_status_prv3;
  assign io_requestor_0_status_fs = io_dpath_status_fs;
  assign io_requestor_0_status_xs = io_dpath_status_xs;
  assign io_requestor_0_status_mprv = io_dpath_status_mprv;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_0_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_0_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_0_status_sd = io_dpath_status_sd;
  assign io_requestor_0_resp_bits_pte_v = r_pte_v;
  assign T210 = T106 ? T71 : r_pte_v;
  assign io_requestor_0_resp_bits_pte_typ = r_pte_typ;
  assign T211 = T106 ? T70 : r_pte_typ;
  assign io_requestor_0_resp_bits_pte_r = r_pte_r;
  assign T212 = T106 ? T114 : r_pte_r;
  assign io_requestor_0_resp_bits_pte_d = r_pte_d;
  assign T213 = T106 ? T111 : r_pte_d;
  assign io_requestor_0_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign T214 = T106 ? T215 : r_pte_reserved_for_software;
  assign T215 = io_mem_resp_bits_data[4'h9:3'h7];
  assign io_requestor_0_resp_bits_pte_ppn = T245;
  assign T245 = resp_ppn[5'h13:1'h0];
  assign resp_ppn = T225 ? r_resp_ppn : T216;
  assign T216 = T223 ? T220 : T217;
  assign T217 = {T219, T218};
  assign T218 = r_req_addr[5'h11:1'h0];
  assign T219 = r_resp_ppn >> 5'h12;
  assign T220 = {T222, T221};
  assign T221 = r_req_addr[4'h8:1'h0];
  assign T222 = r_resp_ppn >> 4'h9;
  assign T223 = T224[1'h0:1'h0];
  assign T224 = count;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hc;
  assign T225 = T224[1'h1:1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = state == 3'h6;
  assign io_requestor_0_resp_valid = T226;
  assign T226 = resp_val & T227;
  assign T227 = r_req_dest == 1'h0;
  assign T228 = T93 ? arb_io_chosen : r_req_dest;
  assign resp_val = T229 | resp_err;
  assign T229 = state == 3'h5;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_ie = io_dpath_status_ie;
  assign io_requestor_1_status_prv = io_dpath_status_prv;
  assign io_requestor_1_status_ie1 = io_dpath_status_ie1;
  assign io_requestor_1_status_prv1 = io_dpath_status_prv1;
  assign io_requestor_1_status_ie2 = io_dpath_status_ie2;
  assign io_requestor_1_status_prv2 = io_dpath_status_prv2;
  assign io_requestor_1_status_ie3 = io_dpath_status_ie3;
  assign io_requestor_1_status_prv3 = io_dpath_status_prv3;
  assign io_requestor_1_status_fs = io_dpath_status_fs;
  assign io_requestor_1_status_xs = io_dpath_status_xs;
  assign io_requestor_1_status_mprv = io_dpath_status_mprv;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_1_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_1_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_1_status_sd = io_dpath_status_sd;
  assign io_requestor_1_resp_bits_pte_v = r_pte_v;
  assign io_requestor_1_resp_bits_pte_typ = r_pte_typ;
  assign io_requestor_1_resp_bits_pte_r = r_pte_r;
  assign io_requestor_1_resp_bits_pte_d = r_pte_d;
  assign io_requestor_1_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_1_resp_bits_pte_ppn = T246;
  assign T246 = resp_ppn[5'h13:1'h0];
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T230;
  assign T230 = resp_val & T231;
  assign T231 = r_req_dest == 1'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  RRArbiter_2 arb(.clk(clk), .reset(reset),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits_addr( io_requestor_1_req_bits_addr ),
       .io_in_1_bits_prv( io_requestor_1_req_bits_prv ),
       .io_in_1_bits_store( io_requestor_1_req_bits_store ),
       .io_in_1_bits_fetch( io_requestor_1_req_bits_fetch ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits_addr( io_requestor_0_req_bits_addr ),
       .io_in_0_bits_prv( io_requestor_0_req_bits_prv ),
       .io_in_0_bits_store( io_requestor_0_req_bits_store ),
       .io_in_0_bits_fetch( io_requestor_0_req_bits_fetch ),
       .io_out_ready( T0 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits_addr( arb_io_out_bits_addr ),
       .io_out_bits_prv( arb_io_out_bits_prv ),
       .io_out_bits_store( arb_io_out_bits_store ),
       .io_out_bits_fetch( arb_io_out_bits_fetch ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T197) begin
      state <= 3'h0;
    end else if(T196) begin
      state <= 3'h0;
    end else if(T195) begin
      state <= 3'h1;
    end else if(T193) begin
      state <= 3'h3;
    end else if(T191) begin
      state <= 3'h4;
    end else if(T188) begin
      state <= T187;
    end else if(T182) begin
      state <= 3'h1;
    end else if(T181) begin
      state <= 3'h6;
    end else if(T179) begin
      state <= 3'h1;
    end else if(T176) begin
      state <= 3'h2;
    end else if(T15) begin
      state <= 3'h1;
    end else if(T13) begin
      state <= 3'h1;
    end
    if(T182) begin
      count <= T22;
    end else if(T15) begin
      count <= T21;
    end else if(T14) begin
      count <= 2'h0;
    end
    if(T72) begin
      R27 <= 1'h0;
    end else if(T30) begin
      R27 <= 1'h1;
    end
    if(T60) begin
      R45 <= T47;
    end
    if(T72) begin
      R73 <= 1'h0;
    end else if(T76) begin
      R73 <= 1'h1;
    end
    if(T72) begin
      R78 <= 1'h0;
    end else if(T81) begin
      R78 <= 1'h1;
    end
    if(T93) begin
      r_req_addr <= arb_io_out_bits_addr;
    end
    if(T15) begin
      r_pte_ppn <= pte_cache_data;
    end else if(T106) begin
      r_pte_ppn <= T105;
    end else if(T93) begin
      r_pte_ppn <= T104;
    end
    if(T93) begin
      r_req_store <= arb_io_out_bits_store;
    end
    if(T93) begin
      r_req_fetch <= arb_io_out_bits_fetch;
    end
    if(T93) begin
      r_req_prv <= arb_io_out_bits_prv;
    end
    if (T154)
      T152[T34] <= T105;
    if (T168)
      T166[T34] <= pte_addr;
    if(T106) begin
      r_pte_v <= T71;
    end
    if(T106) begin
      r_pte_typ <= T70;
    end
    if(T106) begin
      r_pte_r <= T114;
    end
    if(T106) begin
      r_pte_d <= T111;
    end
    if(T106) begin
      r_pte_reserved_for_software <= T215;
    end
    if(T93) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [39:0] io_requestor_1_req_bits_addr,
    input [8:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    input [2:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_kill,
    input  io_requestor_1_req_bits_phys,
    input [63:0] io_requestor_1_req_bits_data,
    output io_requestor_1_resp_valid,
    output[39:0] io_requestor_1_resp_bits_addr,
    output[8:0] io_requestor_1_resp_bits_tag,
    output[4:0] io_requestor_1_resp_bits_cmd,
    output[2:0] io_requestor_1_resp_bits_typ,
    output[63:0] io_requestor_1_resp_bits_data,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data_word_bypass,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[8:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    input  io_requestor_1_invalidate_lr,
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [39:0] io_requestor_0_req_bits_addr,
    input [8:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    input [2:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_kill,
    input  io_requestor_0_req_bits_phys,
    input [63:0] io_requestor_0_req_bits_data,
    output io_requestor_0_resp_valid,
    output[39:0] io_requestor_0_resp_bits_addr,
    output[8:0] io_requestor_0_resp_bits_tag,
    output[4:0] io_requestor_0_resp_bits_cmd,
    output[2:0] io_requestor_0_resp_bits_typ,
    output[63:0] io_requestor_0_resp_bits_data,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data_word_bypass,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[8:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_invalidate_lr
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[39:0] io_mem_req_bits_addr,
    output[8:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_kill,
    output io_mem_req_bits_phys,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [39:0] io_mem_resp_bits_addr,
    input [8:0] io_mem_resp_bits_tag,
    input [4:0] io_mem_resp_bits_cmd,
    input [2:0] io_mem_resp_bits_typ,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_word_bypass,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [8:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_invalidate_lr
    input  io_mem_ordered
);

  wire[63:0] T0;
  reg  r_valid_0;
  wire T1;
  wire T2;
  wire[2:0] T3;
  wire[4:0] T4;
  wire[8:0] T32;
  wire[9:0] T5;
  wire[9:0] T6;
  wire[9:0] T7;
  wire[39:0] T8;
  wire T9;
  wire[8:0] T33;
  wire[7:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[8:0] T34;
  wire[7:0] T18;
  wire T19;
  wire[8:0] T35;
  wire[7:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[8:0] T36;
  wire[7:0] T28;
  wire T29;
  wire T30;
  wire T31;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_valid_0 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_invalidate_lr = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_req_bits_data = T0;
  assign T0 = r_valid_0 ? io_requestor_0_req_bits_data : io_requestor_1_req_bits_data;
  assign io_mem_req_bits_phys = T1;
  assign T1 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign io_mem_req_bits_kill = T2;
  assign T2 = r_valid_0 ? io_requestor_0_req_bits_kill : io_requestor_1_req_bits_kill;
  assign io_mem_req_bits_typ = T3;
  assign T3 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign io_mem_req_bits_cmd = T4;
  assign T4 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign io_mem_req_bits_tag = T32;
  assign T32 = T5[4'h8:1'h0];
  assign T5 = io_requestor_0_req_valid ? T7 : T6;
  assign T6 = {io_requestor_1_req_bits_tag, 1'h1};
  assign T7 = {io_requestor_0_req_bits_tag, 1'h0};
  assign io_mem_req_bits_addr = T8;
  assign T8 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign io_mem_req_valid = T9;
  assign T9 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T33;
  assign T33 = {1'h0, T10};
  assign T10 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_0_replay_next_valid = T11;
  assign T11 = io_mem_replay_next_valid & T12;
  assign T12 = T13 == 1'h0;
  assign T13 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_replay = T14;
  assign T14 = io_mem_resp_bits_replay & T15;
  assign T15 = T16 == 1'h0;
  assign T16 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_0_resp_bits_nack = T17;
  assign T17 = io_mem_resp_bits_nack & T15;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T34;
  assign T34 = {1'h0, T18};
  assign T18 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_valid = T19;
  assign T19 = io_mem_resp_valid & T15;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T35;
  assign T35 = {1'h0, T20};
  assign T20 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_1_replay_next_valid = T21;
  assign T21 = io_mem_replay_next_valid & T22;
  assign T22 = T23 == 1'h1;
  assign T23 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_replay = T24;
  assign T24 = io_mem_resp_bits_replay & T25;
  assign T25 = T26 == 1'h1;
  assign T26 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_1_resp_bits_nack = T27;
  assign T27 = io_mem_resp_bits_nack & T25;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T36;
  assign T36 = {1'h0, T28};
  assign T28 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_valid = T29;
  assign T29 = io_mem_resp_valid & T25;
  assign io_requestor_1_req_ready = T30;
  assign T30 = io_requestor_0_req_ready & T31;
  assign T31 = io_requestor_0_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module RocketTile(input clk, input reset,
    input  io_cached_0_acquire_ready,
    output io_cached_0_acquire_valid,
    output[25:0] io_cached_0_acquire_bits_addr_block,
    output[1:0] io_cached_0_acquire_bits_client_xact_id,
    output[1:0] io_cached_0_acquire_bits_addr_beat,
    output io_cached_0_acquire_bits_is_builtin_type,
    output[2:0] io_cached_0_acquire_bits_a_type,
    output[16:0] io_cached_0_acquire_bits_union,
    output[127:0] io_cached_0_acquire_bits_data,
    output io_cached_0_grant_ready,
    input  io_cached_0_grant_valid,
    input [1:0] io_cached_0_grant_bits_addr_beat,
    input [1:0] io_cached_0_grant_bits_client_xact_id,
    input [3:0] io_cached_0_grant_bits_manager_xact_id,
    input  io_cached_0_grant_bits_is_builtin_type,
    input [3:0] io_cached_0_grant_bits_g_type,
    input [127:0] io_cached_0_grant_bits_data,
    output io_cached_0_probe_ready,
    input  io_cached_0_probe_valid,
    input [25:0] io_cached_0_probe_bits_addr_block,
    input [1:0] io_cached_0_probe_bits_p_type,
    input  io_cached_0_release_ready,
    output io_cached_0_release_valid,
    output[1:0] io_cached_0_release_bits_addr_beat,
    output[25:0] io_cached_0_release_bits_addr_block,
    output[1:0] io_cached_0_release_bits_client_xact_id,
    output[2:0] io_cached_0_release_bits_r_type,
    output io_cached_0_release_bits_voluntary,
    output[127:0] io_cached_0_release_bits_data,
    input  io_uncached_0_acquire_ready,
    output io_uncached_0_acquire_valid,
    output[25:0] io_uncached_0_acquire_bits_addr_block,
    output[1:0] io_uncached_0_acquire_bits_client_xact_id,
    output[1:0] io_uncached_0_acquire_bits_addr_beat,
    output io_uncached_0_acquire_bits_is_builtin_type,
    output[2:0] io_uncached_0_acquire_bits_a_type,
    output[16:0] io_uncached_0_acquire_bits_union,
    output[127:0] io_uncached_0_acquire_bits_data,
    output io_uncached_0_grant_ready,
    input  io_uncached_0_grant_valid,
    input [1:0] io_uncached_0_grant_bits_addr_beat,
    input [1:0] io_uncached_0_grant_bits_client_xact_id,
    input [3:0] io_uncached_0_grant_bits_manager_xact_id,
    input  io_uncached_0_grant_bits_is_builtin_type,
    input [3:0] io_uncached_0_grant_bits_g_type,
    input [127:0] io_uncached_0_grant_bits_data,
    input  io_host_reset,
    input  io_host_id,
    output io_host_csr_req_ready,
    input  io_host_csr_req_valid,
    input  io_host_csr_req_bits_rw,
    input [11:0] io_host_csr_req_bits_addr,
    input [63:0] io_host_csr_req_bits_data,
    input  io_host_csr_resp_ready,
    output io_host_csr_resp_valid,
    output[63:0] io_host_csr_resp_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_csr
);

  wire dcArb_io_requestor_1_req_ready;
  wire dcArb_io_requestor_1_resp_valid;
  wire[39:0] dcArb_io_requestor_1_resp_bits_addr;
  wire[8:0] dcArb_io_requestor_1_resp_bits_tag;
  wire[4:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire[2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data;
  wire dcArb_io_requestor_1_resp_bits_nack;
  wire dcArb_io_requestor_1_resp_bits_replay;
  wire dcArb_io_requestor_1_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data_word_bypass;
  wire[63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire dcArb_io_requestor_1_replay_next_valid;
  wire[8:0] dcArb_io_requestor_1_replay_next_bits;
  wire dcArb_io_requestor_1_xcpt_ma_ld;
  wire dcArb_io_requestor_1_xcpt_ma_st;
  wire dcArb_io_requestor_1_xcpt_pf_ld;
  wire dcArb_io_requestor_1_xcpt_pf_st;
  wire dcArb_io_requestor_1_ordered;
  wire dcArb_io_requestor_0_req_ready;
  wire dcArb_io_requestor_0_resp_valid;
  wire[39:0] dcArb_io_requestor_0_resp_bits_addr;
  wire[8:0] dcArb_io_requestor_0_resp_bits_tag;
  wire[4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire[2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data;
  wire dcArb_io_requestor_0_resp_bits_nack;
  wire dcArb_io_requestor_0_resp_bits_replay;
  wire dcArb_io_requestor_0_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data_word_bypass;
  wire[63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire dcArb_io_requestor_0_replay_next_valid;
  wire[8:0] dcArb_io_requestor_0_replay_next_bits;
  wire dcArb_io_requestor_0_xcpt_ma_ld;
  wire dcArb_io_requestor_0_xcpt_ma_st;
  wire dcArb_io_requestor_0_xcpt_pf_ld;
  wire dcArb_io_requestor_0_xcpt_pf_st;
  wire dcArb_io_requestor_0_ordered;
  wire dcArb_io_mem_req_valid;
  wire[39:0] dcArb_io_mem_req_bits_addr;
  wire[8:0] dcArb_io_mem_req_bits_tag;
  wire[4:0] dcArb_io_mem_req_bits_cmd;
  wire[2:0] dcArb_io_mem_req_bits_typ;
  wire dcArb_io_mem_req_bits_kill;
  wire dcArb_io_mem_req_bits_phys;
  wire[63:0] dcArb_io_mem_req_bits_data;
  wire core_io_host_csr_req_ready;
  wire core_io_host_csr_resp_valid;
  wire[63:0] core_io_host_csr_resp_bits;
  wire core_io_host_ipi_req_valid;
  wire core_io_host_ipi_req_bits;
  wire core_io_host_ipi_rep_ready;
  wire core_io_host_debug_stats_csr;
  wire core_io_imem_req_valid;
  wire[39:0] core_io_imem_req_bits_pc;
  wire core_io_imem_resp_ready;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire core_io_imem_btb_update_bits_prediction_bits_mask;
  wire core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[38:0] core_io_imem_btb_update_bits_pc;
  wire[38:0] core_io_imem_btb_update_bits_target;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_isReturn;
  wire[38:0] core_io_imem_btb_update_bits_br_pc;
  wire core_io_imem_bht_update_valid;
  wire core_io_imem_bht_update_bits_prediction_valid;
  wire core_io_imem_bht_update_bits_prediction_bits_taken;
  wire core_io_imem_bht_update_bits_prediction_bits_mask;
  wire core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_bht_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire[38:0] core_io_imem_bht_update_bits_pc;
  wire core_io_imem_bht_update_bits_taken;
  wire core_io_imem_bht_update_bits_mispredict;
  wire core_io_imem_ras_update_valid;
  wire core_io_imem_ras_update_bits_isCall;
  wire core_io_imem_ras_update_bits_isReturn;
  wire[38:0] core_io_imem_ras_update_bits_returnAddr;
  wire core_io_imem_ras_update_bits_prediction_valid;
  wire core_io_imem_ras_update_bits_prediction_bits_taken;
  wire core_io_imem_ras_update_bits_prediction_bits_mask;
  wire core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_ras_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire core_io_imem_invalidate;
  wire core_io_dmem_req_valid;
  wire[39:0] core_io_dmem_req_bits_addr;
  wire[8:0] core_io_dmem_req_bits_tag;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[2:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_kill;
  wire core_io_dmem_req_bits_phys;
  wire[63:0] core_io_dmem_req_bits_data;
  wire core_io_dmem_invalidate_lr;
  wire[31:0] core_io_ptw_ptbr;
  wire core_io_ptw_invalidate;
  wire core_io_ptw_status_sd;
  wire[30:0] core_io_ptw_status_zero2;
  wire core_io_ptw_status_sd_rv32;
  wire[8:0] core_io_ptw_status_zero1;
  wire[4:0] core_io_ptw_status_vm;
  wire core_io_ptw_status_mprv;
  wire[1:0] core_io_ptw_status_xs;
  wire[1:0] core_io_ptw_status_fs;
  wire[1:0] core_io_ptw_status_prv3;
  wire core_io_ptw_status_ie3;
  wire[1:0] core_io_ptw_status_prv2;
  wire core_io_ptw_status_ie2;
  wire[1:0] core_io_ptw_status_prv1;
  wire core_io_ptw_status_ie1;
  wire[1:0] core_io_ptw_status_prv;
  wire core_io_ptw_status_ie;
  wire ptw_io_requestor_1_req_ready;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_resp_bits_error;
  wire[19:0] ptw_io_requestor_1_resp_bits_pte_ppn;
  wire[2:0] ptw_io_requestor_1_resp_bits_pte_reserved_for_software;
  wire ptw_io_requestor_1_resp_bits_pte_d;
  wire ptw_io_requestor_1_resp_bits_pte_r;
  wire[3:0] ptw_io_requestor_1_resp_bits_pte_typ;
  wire ptw_io_requestor_1_resp_bits_pte_v;
  wire ptw_io_requestor_1_status_sd;
  wire[30:0] ptw_io_requestor_1_status_zero2;
  wire ptw_io_requestor_1_status_sd_rv32;
  wire[8:0] ptw_io_requestor_1_status_zero1;
  wire[4:0] ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_mprv;
  wire[1:0] ptw_io_requestor_1_status_xs;
  wire[1:0] ptw_io_requestor_1_status_fs;
  wire[1:0] ptw_io_requestor_1_status_prv3;
  wire ptw_io_requestor_1_status_ie3;
  wire[1:0] ptw_io_requestor_1_status_prv2;
  wire ptw_io_requestor_1_status_ie2;
  wire[1:0] ptw_io_requestor_1_status_prv1;
  wire ptw_io_requestor_1_status_ie1;
  wire[1:0] ptw_io_requestor_1_status_prv;
  wire ptw_io_requestor_1_status_ie;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_0_req_ready;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_resp_bits_error;
  wire[19:0] ptw_io_requestor_0_resp_bits_pte_ppn;
  wire[2:0] ptw_io_requestor_0_resp_bits_pte_reserved_for_software;
  wire ptw_io_requestor_0_resp_bits_pte_d;
  wire ptw_io_requestor_0_resp_bits_pte_r;
  wire[3:0] ptw_io_requestor_0_resp_bits_pte_typ;
  wire ptw_io_requestor_0_resp_bits_pte_v;
  wire ptw_io_requestor_0_status_sd;
  wire[30:0] ptw_io_requestor_0_status_zero2;
  wire ptw_io_requestor_0_status_sd_rv32;
  wire[8:0] ptw_io_requestor_0_status_zero1;
  wire[4:0] ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_mprv;
  wire[1:0] ptw_io_requestor_0_status_xs;
  wire[1:0] ptw_io_requestor_0_status_fs;
  wire[1:0] ptw_io_requestor_0_status_prv3;
  wire ptw_io_requestor_0_status_ie3;
  wire[1:0] ptw_io_requestor_0_status_prv2;
  wire ptw_io_requestor_0_status_ie2;
  wire[1:0] ptw_io_requestor_0_status_prv1;
  wire ptw_io_requestor_0_status_ie1;
  wire[1:0] ptw_io_requestor_0_status_prv;
  wire ptw_io_requestor_0_status_ie;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_mem_req_valid;
  wire[39:0] ptw_io_mem_req_bits_addr;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire[2:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_kill;
  wire ptw_io_mem_req_bits_phys;
  wire[63:0] ptw_io_mem_req_bits_data;
  wire icache_io_cpu_resp_valid;
  wire[39:0] icache_io_cpu_resp_bits_pc;
  wire[31:0] icache_io_cpu_resp_bits_data_0;
  wire icache_io_cpu_resp_bits_mask;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire icache_io_cpu_btb_resp_bits_mask;
  wire icache_io_cpu_btb_resp_bits_bridx;
  wire[38:0] icache_io_cpu_btb_resp_bits_target;
  wire[5:0] icache_io_cpu_btb_resp_bits_entry;
  wire[6:0] icache_io_cpu_btb_resp_bits_bht_history;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire[39:0] icache_io_cpu_npc;
  wire icache_io_ptw_req_valid;
  wire[26:0] icache_io_ptw_req_bits_addr;
  wire[1:0] icache_io_ptw_req_bits_prv;
  wire icache_io_ptw_req_bits_store;
  wire icache_io_ptw_req_bits_fetch;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_addr_block;
  wire[1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] icache_io_mem_acquire_bits_addr_beat;
  wire icache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] icache_io_mem_acquire_bits_a_type;
  wire[16:0] icache_io_mem_acquire_bits_union;
  wire[127:0] icache_io_mem_acquire_bits_data;
  wire icache_io_mem_grant_ready;
  wire dcache_io_cpu_req_ready;
  wire dcache_io_cpu_resp_valid;
  wire[39:0] dcache_io_cpu_resp_bits_addr;
  wire[8:0] dcache_io_cpu_resp_bits_tag;
  wire[4:0] dcache_io_cpu_resp_bits_cmd;
  wire[2:0] dcache_io_cpu_resp_bits_typ;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_bits_replay;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[63:0] dcache_io_cpu_resp_bits_data_word_bypass;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire dcache_io_cpu_replay_next_valid;
  wire[8:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_ordered;
  wire dcache_io_ptw_req_valid;
  wire[26:0] dcache_io_ptw_req_bits_addr;
  wire[1:0] dcache_io_ptw_req_bits_prv;
  wire dcache_io_ptw_req_bits_store;
  wire dcache_io_ptw_req_bits_fetch;
  wire dcache_io_mem_acquire_valid;
  wire[25:0] dcache_io_mem_acquire_bits_addr_block;
  wire[1:0] dcache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] dcache_io_mem_acquire_bits_addr_beat;
  wire dcache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] dcache_io_mem_acquire_bits_a_type;
  wire[16:0] dcache_io_mem_acquire_bits_union;
  wire[127:0] dcache_io_mem_acquire_bits_data;
  wire dcache_io_mem_grant_ready;
  wire dcache_io_mem_probe_ready;
  wire dcache_io_mem_release_valid;
  wire[1:0] dcache_io_mem_release_bits_addr_beat;
  wire[25:0] dcache_io_mem_release_bits_addr_block;
  wire[1:0] dcache_io_mem_release_bits_client_xact_id;
  wire[2:0] dcache_io_mem_release_bits_r_type;
  wire dcache_io_mem_release_bits_voluntary;
  wire[127:0] dcache_io_mem_release_bits_data;


  assign io_host_debug_stats_csr = core_io_host_debug_stats_csr;
  assign io_host_ipi_rep_ready = core_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = core_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = core_io_host_ipi_req_valid;
  assign io_host_csr_resp_bits = core_io_host_csr_resp_bits;
  assign io_host_csr_resp_valid = core_io_host_csr_resp_valid;
  assign io_host_csr_req_ready = core_io_host_csr_req_ready;
  assign io_uncached_0_grant_ready = icache_io_mem_grant_ready;
  assign io_uncached_0_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_uncached_0_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_uncached_0_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_uncached_0_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_uncached_0_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_uncached_0_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_uncached_0_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_uncached_0_acquire_valid = icache_io_mem_acquire_valid;
  assign io_cached_0_release_bits_data = dcache_io_mem_release_bits_data;
  assign io_cached_0_release_bits_voluntary = dcache_io_mem_release_bits_voluntary;
  assign io_cached_0_release_bits_r_type = dcache_io_mem_release_bits_r_type;
  assign io_cached_0_release_bits_client_xact_id = dcache_io_mem_release_bits_client_xact_id;
  assign io_cached_0_release_bits_addr_block = dcache_io_mem_release_bits_addr_block;
  assign io_cached_0_release_bits_addr_beat = dcache_io_mem_release_bits_addr_beat;
  assign io_cached_0_release_valid = dcache_io_mem_release_valid;
  assign io_cached_0_probe_ready = dcache_io_mem_probe_ready;
  assign io_cached_0_grant_ready = dcache_io_mem_grant_ready;
  assign io_cached_0_acquire_bits_data = dcache_io_mem_acquire_bits_data;
  assign io_cached_0_acquire_bits_union = dcache_io_mem_acquire_bits_union;
  assign io_cached_0_acquire_bits_a_type = dcache_io_mem_acquire_bits_a_type;
  assign io_cached_0_acquire_bits_is_builtin_type = dcache_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_0_acquire_bits_addr_beat = dcache_io_mem_acquire_bits_addr_beat;
  assign io_cached_0_acquire_bits_client_xact_id = dcache_io_mem_acquire_bits_client_xact_id;
  assign io_cached_0_acquire_bits_addr_block = dcache_io_mem_acquire_bits_addr_block;
  assign io_cached_0_acquire_valid = dcache_io_mem_acquire_valid;
  Rocket core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_csr_req_ready( core_io_host_csr_req_ready ),
       .io_host_csr_req_valid( io_host_csr_req_valid ),
       .io_host_csr_req_bits_rw( io_host_csr_req_bits_rw ),
       .io_host_csr_req_bits_addr( io_host_csr_req_bits_addr ),
       .io_host_csr_req_bits_data( io_host_csr_req_bits_data ),
       .io_host_csr_resp_ready( io_host_csr_resp_ready ),
       .io_host_csr_resp_valid( core_io_host_csr_resp_valid ),
       .io_host_csr_resp_bits( core_io_host_csr_resp_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( core_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( core_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( core_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_csr( core_io_host_debug_stats_csr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_imem_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_imem_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_imem_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_imem_btb_update_bits_taken(  )
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_imem_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_imem_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_imem_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_imem_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_imem_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_imem_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_imem_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_imem_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_imem_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_imem_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_imem_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_imem_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_imem_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_imem_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_imem_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_imem_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_imem_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_imem_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_imem_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_imem_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_imem_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_imem_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_imem_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_imem_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_imem_npc( icache_io_cpu_npc ),
       .io_dmem_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data_word_bypass( dcArb_io_requestor_1_resp_bits_data_word_bypass ),
       .io_dmem_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       .io_dmem_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_dmem_ordered( dcArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_status_sd( core_io_ptw_status_sd ),
       .io_ptw_status_zero2( core_io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( core_io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( core_io_ptw_status_zero1 ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_mprv( core_io_ptw_status_mprv ),
       .io_ptw_status_xs( core_io_ptw_status_xs ),
       .io_ptw_status_fs( core_io_ptw_status_fs ),
       .io_ptw_status_prv3( core_io_ptw_status_prv3 ),
       .io_ptw_status_ie3( core_io_ptw_status_ie3 ),
       .io_ptw_status_prv2( core_io_ptw_status_prv2 ),
       .io_ptw_status_ie2( core_io_ptw_status_ie2 ),
       .io_ptw_status_prv1( core_io_ptw_status_prv1 ),
       .io_ptw_status_ie1( core_io_ptw_status_ie1 ),
       .io_ptw_status_prv( core_io_ptw_status_prv ),
       .io_ptw_status_ie( core_io_ptw_status_ie )
       //.io_fpu_inst(  )
       //.io_fpu_fromint_data(  )
       //.io_fpu_fcsr_rm(  )
       //.io_fpu_fcsr_flags_valid(  )
       //.io_fpu_fcsr_flags_bits(  )
       //.io_fpu_store_data(  )
       //.io_fpu_toint_data(  )
       //.io_fpu_dmem_resp_val(  )
       //.io_fpu_dmem_resp_type(  )
       //.io_fpu_dmem_resp_tag(  )
       //.io_fpu_dmem_resp_data(  )
       //.io_fpu_valid(  )
       //.io_fpu_fcsr_rdy(  )
       //.io_fpu_nack_mem(  )
       //.io_fpu_illegal_rm(  )
       //.io_fpu_killx(  )
       //.io_fpu_killm(  )
       //.io_fpu_dec_cmd(  )
       //.io_fpu_dec_ldst(  )
       //.io_fpu_dec_wen(  )
       //.io_fpu_dec_ren1(  )
       //.io_fpu_dec_ren2(  )
       //.io_fpu_dec_ren3(  )
       //.io_fpu_dec_swap12(  )
       //.io_fpu_dec_swap23(  )
       //.io_fpu_dec_single(  )
       //.io_fpu_dec_fromint(  )
       //.io_fpu_dec_toint(  )
       //.io_fpu_dec_fastpipe(  )
       //.io_fpu_dec_fma(  )
       //.io_fpu_dec_div(  )
       //.io_fpu_dec_sqrt(  )
       //.io_fpu_dec_round(  )
       //.io_fpu_dec_wflags(  )
       //.io_fpu_sboard_set(  )
       //.io_fpu_sboard_clr(  )
       //.io_fpu_sboard_clra(  )
       //.io_rocc_cmd_ready(  )
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       //.io_rocc_resp_valid(  )
       //.io_rocc_resp_bits_rd(  )
       //.io_rocc_resp_bits_data(  )
       //.io_rocc_mem_req_ready(  )
       //.io_rocc_mem_req_valid(  )
       //.io_rocc_mem_req_bits_addr(  )
       //.io_rocc_mem_req_bits_tag(  )
       //.io_rocc_mem_req_bits_cmd(  )
       //.io_rocc_mem_req_bits_typ(  )
       //.io_rocc_mem_req_bits_kill(  )
       //.io_rocc_mem_req_bits_phys(  )
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_word_bypass(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_invalidate_lr(  )
       //.io_rocc_mem_ordered(  )
       //.io_rocc_busy(  )
       //.io_rocc_s(  )
       //.io_rocc_interrupt(  )
       //.io_rocc_imem_acquire_ready(  )
       //.io_rocc_imem_acquire_valid(  )
       //.io_rocc_imem_acquire_bits_addr_block(  )
       //.io_rocc_imem_acquire_bits_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_addr_beat(  )
       //.io_rocc_imem_acquire_bits_is_builtin_type(  )
       //.io_rocc_imem_acquire_bits_a_type(  )
       //.io_rocc_imem_acquire_bits_union(  )
       //.io_rocc_imem_acquire_bits_data(  )
       //.io_rocc_imem_grant_ready(  )
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_addr_beat(  )
       //.io_rocc_imem_grant_bits_client_xact_id(  )
       //.io_rocc_imem_grant_bits_manager_xact_id(  )
       //.io_rocc_imem_grant_bits_is_builtin_type(  )
       //.io_rocc_imem_grant_bits_g_type(  )
       //.io_rocc_imem_grant_bits_data(  )
       //.io_rocc_dmem_0_acquire_ready(  )
       //.io_rocc_dmem_0_acquire_valid(  )
       //.io_rocc_dmem_0_acquire_bits_addr_block(  )
       //.io_rocc_dmem_0_acquire_bits_client_xact_id(  )
       //.io_rocc_dmem_0_acquire_bits_addr_beat(  )
       //.io_rocc_dmem_0_acquire_bits_is_builtin_type(  )
       //.io_rocc_dmem_0_acquire_bits_a_type(  )
       //.io_rocc_dmem_0_acquire_bits_union(  )
       //.io_rocc_dmem_0_acquire_bits_data(  )
       //.io_rocc_dmem_0_grant_ready(  )
       //.io_rocc_dmem_0_grant_valid(  )
       //.io_rocc_dmem_0_grant_bits_addr_beat(  )
       //.io_rocc_dmem_0_grant_bits_client_xact_id(  )
       //.io_rocc_dmem_0_grant_bits_manager_xact_id(  )
       //.io_rocc_dmem_0_grant_bits_is_builtin_type(  )
       //.io_rocc_dmem_0_grant_bits_g_type(  )
       //.io_rocc_dmem_0_grant_bits_data(  )
       //.io_rocc_iptw_req_ready(  )
       //.io_rocc_iptw_req_valid(  )
       //.io_rocc_iptw_req_bits_addr(  )
       //.io_rocc_iptw_req_bits_prv(  )
       //.io_rocc_iptw_req_bits_store(  )
       //.io_rocc_iptw_req_bits_fetch(  )
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_pte_ppn(  )
       //.io_rocc_iptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_iptw_resp_bits_pte_d(  )
       //.io_rocc_iptw_resp_bits_pte_r(  )
       //.io_rocc_iptw_resp_bits_pte_typ(  )
       //.io_rocc_iptw_resp_bits_pte_v(  )
       //.io_rocc_iptw_status_sd(  )
       //.io_rocc_iptw_status_zero2(  )
       //.io_rocc_iptw_status_sd_rv32(  )
       //.io_rocc_iptw_status_zero1(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_mprv(  )
       //.io_rocc_iptw_status_xs(  )
       //.io_rocc_iptw_status_fs(  )
       //.io_rocc_iptw_status_prv3(  )
       //.io_rocc_iptw_status_ie3(  )
       //.io_rocc_iptw_status_prv2(  )
       //.io_rocc_iptw_status_ie2(  )
       //.io_rocc_iptw_status_prv1(  )
       //.io_rocc_iptw_status_ie1(  )
       //.io_rocc_iptw_status_prv(  )
       //.io_rocc_iptw_status_ie(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_dptw_req_ready(  )
       //.io_rocc_dptw_req_valid(  )
       //.io_rocc_dptw_req_bits_addr(  )
       //.io_rocc_dptw_req_bits_prv(  )
       //.io_rocc_dptw_req_bits_store(  )
       //.io_rocc_dptw_req_bits_fetch(  )
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_pte_ppn(  )
       //.io_rocc_dptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_dptw_resp_bits_pte_d(  )
       //.io_rocc_dptw_resp_bits_pte_r(  )
       //.io_rocc_dptw_resp_bits_pte_typ(  )
       //.io_rocc_dptw_resp_bits_pte_v(  )
       //.io_rocc_dptw_status_sd(  )
       //.io_rocc_dptw_status_zero2(  )
       //.io_rocc_dptw_status_sd_rv32(  )
       //.io_rocc_dptw_status_zero1(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_mprv(  )
       //.io_rocc_dptw_status_xs(  )
       //.io_rocc_dptw_status_fs(  )
       //.io_rocc_dptw_status_prv3(  )
       //.io_rocc_dptw_status_ie3(  )
       //.io_rocc_dptw_status_prv2(  )
       //.io_rocc_dptw_status_ie2(  )
       //.io_rocc_dptw_status_prv1(  )
       //.io_rocc_dptw_status_ie1(  )
       //.io_rocc_dptw_status_prv(  )
       //.io_rocc_dptw_status_ie(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_pptw_req_ready(  )
       //.io_rocc_pptw_req_valid(  )
       //.io_rocc_pptw_req_bits_addr(  )
       //.io_rocc_pptw_req_bits_prv(  )
       //.io_rocc_pptw_req_bits_store(  )
       //.io_rocc_pptw_req_bits_fetch(  )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_pte_ppn(  )
       //.io_rocc_pptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_pptw_resp_bits_pte_d(  )
       //.io_rocc_pptw_resp_bits_pte_r(  )
       //.io_rocc_pptw_resp_bits_pte_typ(  )
       //.io_rocc_pptw_resp_bits_pte_v(  )
       //.io_rocc_pptw_status_sd(  )
       //.io_rocc_pptw_status_zero2(  )
       //.io_rocc_pptw_status_sd_rv32(  )
       //.io_rocc_pptw_status_zero1(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_mprv(  )
       //.io_rocc_pptw_status_xs(  )
       //.io_rocc_pptw_status_fs(  )
       //.io_rocc_pptw_status_prv3(  )
       //.io_rocc_pptw_status_ie3(  )
       //.io_rocc_pptw_status_prv2(  )
       //.io_rocc_pptw_status_ie2(  )
       //.io_rocc_pptw_status_prv1(  )
       //.io_rocc_pptw_status_ie1(  )
       //.io_rocc_pptw_status_prv(  )
       //.io_rocc_pptw_status_ie(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_exception(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign core.io_fpu_fcsr_flags_valid = {1{$random}};
    assign core.io_fpu_fcsr_flags_bits = {1{$random}};
    assign core.io_fpu_store_data = {2{$random}};
    assign core.io_fpu_toint_data = {2{$random}};
    assign core.io_fpu_nack_mem = {1{$random}};
    assign core.io_fpu_illegal_rm = {1{$random}};
    assign core.io_fpu_dec_wen = {1{$random}};
    assign core.io_fpu_dec_ren1 = {1{$random}};
    assign core.io_fpu_dec_ren2 = {1{$random}};
    assign core.io_fpu_dec_ren3 = {1{$random}};
    assign core.io_rocc_cmd_ready = {1{$random}};
    assign core.io_rocc_resp_valid = {1{$random}};
    assign core.io_rocc_resp_bits_rd = {1{$random}};
    assign core.io_rocc_resp_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_valid = {1{$random}};
    assign core.io_rocc_mem_req_bits_addr = {2{$random}};
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_cmd = {1{$random}};
    assign core.io_rocc_mem_req_bits_typ = {1{$random}};
    assign core.io_rocc_mem_req_bits_kill = {1{$random}};
    assign core.io_rocc_mem_req_bits_phys = {1{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_invalidate_lr = {1{$random}};
    assign core.io_rocc_busy = {1{$random}};
    assign core.io_rocc_interrupt = {1{$random}};
    assign core.io_rocc_imem_acquire_valid = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_addr_block = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_client_xact_id = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_addr_beat = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_is_builtin_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_a_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_union = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_data = {4{$random}};
    assign core.io_rocc_imem_grant_ready = {1{$random}};
    assign core.io_rocc_dmem_0_acquire_valid = {1{$random}};
    assign core.io_rocc_dmem_0_acquire_bits_addr_block = {1{$random}};
    assign core.io_rocc_dmem_0_acquire_bits_client_xact_id = {1{$random}};
    assign core.io_rocc_dmem_0_acquire_bits_addr_beat = {1{$random}};
    assign core.io_rocc_dmem_0_acquire_bits_is_builtin_type = {1{$random}};
    assign core.io_rocc_dmem_0_acquire_bits_a_type = {1{$random}};
    assign core.io_rocc_dmem_0_acquire_bits_union = {1{$random}};
    assign core.io_rocc_dmem_0_acquire_bits_data = {4{$random}};
    assign core.io_rocc_dmem_0_grant_ready = {1{$random}};
    assign core.io_rocc_iptw_req_valid = {1{$random}};
    assign core.io_rocc_iptw_req_bits_addr = {1{$random}};
    assign core.io_rocc_iptw_req_bits_prv = {1{$random}};
    assign core.io_rocc_iptw_req_bits_store = {1{$random}};
    assign core.io_rocc_iptw_req_bits_fetch = {1{$random}};
    assign core.io_rocc_dptw_req_valid = {1{$random}};
    assign core.io_rocc_dptw_req_bits_addr = {1{$random}};
    assign core.io_rocc_dptw_req_bits_prv = {1{$random}};
    assign core.io_rocc_dptw_req_bits_store = {1{$random}};
    assign core.io_rocc_dptw_req_bits_fetch = {1{$random}};
    assign core.io_rocc_pptw_req_valid = {1{$random}};
    assign core.io_rocc_pptw_req_bits_addr = {1{$random}};
    assign core.io_rocc_pptw_req_bits_prv = {1{$random}};
    assign core.io_rocc_pptw_req_bits_store = {1{$random}};
    assign core.io_rocc_pptw_req_bits_fetch = {1{$random}};
// synthesis translate_on
`endif
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_cpu_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_cpu_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_cpu_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_cpu_btb_update_bits_taken(  )
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_cpu_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_cpu_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_cpu_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_cpu_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_cpu_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_cpu_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_cpu_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_cpu_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_cpu_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_cpu_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_cpu_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_cpu_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_cpu_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_cpu_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_cpu_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_cpu_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_cpu_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_cpu_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_cpu_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_cpu_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_cpu_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_cpu_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_cpu_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_cpu_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_cpu_npc( icache_io_cpu_npc ),
       .io_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_ptw_req_valid( icache_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( icache_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( icache_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( icache_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( icache_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( ptw_io_requestor_0_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( ptw_io_requestor_0_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( ptw_io_requestor_0_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( ptw_io_requestor_0_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( ptw_io_requestor_0_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( ptw_io_requestor_0_resp_bits_pte_v ),
       .io_ptw_status_sd( ptw_io_requestor_0_status_sd ),
       .io_ptw_status_zero2( ptw_io_requestor_0_status_zero2 ),
       .io_ptw_status_sd_rv32( ptw_io_requestor_0_status_sd_rv32 ),
       .io_ptw_status_zero1( ptw_io_requestor_0_status_zero1 ),
       .io_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_ptw_status_mprv( ptw_io_requestor_0_status_mprv ),
       .io_ptw_status_xs( ptw_io_requestor_0_status_xs ),
       .io_ptw_status_fs( ptw_io_requestor_0_status_fs ),
       .io_ptw_status_prv3( ptw_io_requestor_0_status_prv3 ),
       .io_ptw_status_ie3( ptw_io_requestor_0_status_ie3 ),
       .io_ptw_status_prv2( ptw_io_requestor_0_status_prv2 ),
       .io_ptw_status_ie2( ptw_io_requestor_0_status_ie2 ),
       .io_ptw_status_prv1( ptw_io_requestor_0_status_prv1 ),
       .io_ptw_status_ie1( ptw_io_requestor_0_status_ie1 ),
       .io_ptw_status_prv( ptw_io_requestor_0_status_prv ),
       .io_ptw_status_ie( ptw_io_requestor_0_status_ie ),
       .io_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_mem_acquire_ready( io_uncached_0_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( icache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( icache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( icache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( icache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( icache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( icache_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( icache_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_uncached_0_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_uncached_0_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_uncached_0_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_uncached_0_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_uncached_0_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_uncached_0_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_uncached_0_grant_bits_data )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign icache.io_cpu_btb_update_bits_taken = {1{$random}};
// synthesis translate_on
`endif
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcArb_io_mem_req_valid ),
       .io_cpu_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_cpu_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data_word_bypass( dcache_io_cpu_resp_bits_data_word_bypass ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_ptw_req_valid( dcache_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( dcache_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( dcache_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( dcache_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( dcache_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( ptw_io_requestor_1_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( ptw_io_requestor_1_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( ptw_io_requestor_1_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( ptw_io_requestor_1_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( ptw_io_requestor_1_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( ptw_io_requestor_1_resp_bits_pte_v ),
       .io_ptw_status_sd( ptw_io_requestor_1_status_sd ),
       .io_ptw_status_zero2( ptw_io_requestor_1_status_zero2 ),
       .io_ptw_status_sd_rv32( ptw_io_requestor_1_status_sd_rv32 ),
       .io_ptw_status_zero1( ptw_io_requestor_1_status_zero1 ),
       .io_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_ptw_status_mprv( ptw_io_requestor_1_status_mprv ),
       .io_ptw_status_xs( ptw_io_requestor_1_status_xs ),
       .io_ptw_status_fs( ptw_io_requestor_1_status_fs ),
       .io_ptw_status_prv3( ptw_io_requestor_1_status_prv3 ),
       .io_ptw_status_ie3( ptw_io_requestor_1_status_ie3 ),
       .io_ptw_status_prv2( ptw_io_requestor_1_status_prv2 ),
       .io_ptw_status_ie2( ptw_io_requestor_1_status_ie2 ),
       .io_ptw_status_prv1( ptw_io_requestor_1_status_prv1 ),
       .io_ptw_status_ie1( ptw_io_requestor_1_status_ie1 ),
       .io_ptw_status_prv( ptw_io_requestor_1_status_prv ),
       .io_ptw_status_ie( ptw_io_requestor_1_status_ie ),
       .io_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_mem_acquire_ready( io_cached_0_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( dcache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( dcache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( dcache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( dcache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( dcache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( dcache_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( dcache_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_cached_0_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_cached_0_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_cached_0_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_cached_0_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_cached_0_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_cached_0_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_cached_0_grant_bits_data ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( io_cached_0_probe_valid ),
       .io_mem_probe_bits_addr_block( io_cached_0_probe_bits_addr_block ),
       .io_mem_probe_bits_p_type( io_cached_0_probe_bits_p_type ),
       .io_mem_release_ready( io_cached_0_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_addr_beat( dcache_io_mem_release_bits_addr_beat ),
       .io_mem_release_bits_addr_block( dcache_io_mem_release_bits_addr_block ),
       .io_mem_release_bits_client_xact_id( dcache_io_mem_release_bits_client_xact_id ),
       .io_mem_release_bits_r_type( dcache_io_mem_release_bits_r_type ),
       .io_mem_release_bits_voluntary( dcache_io_mem_release_bits_voluntary ),
       .io_mem_release_bits_data( dcache_io_mem_release_bits_data )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_ptw_req_valid ),
       .io_requestor_1_req_bits_addr( dcache_io_ptw_req_bits_addr ),
       .io_requestor_1_req_bits_prv( dcache_io_ptw_req_bits_prv ),
       .io_requestor_1_req_bits_store( dcache_io_ptw_req_bits_store ),
       .io_requestor_1_req_bits_fetch( dcache_io_ptw_req_bits_fetch ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_pte_ppn( ptw_io_requestor_1_resp_bits_pte_ppn ),
       .io_requestor_1_resp_bits_pte_reserved_for_software( ptw_io_requestor_1_resp_bits_pte_reserved_for_software ),
       .io_requestor_1_resp_bits_pte_d( ptw_io_requestor_1_resp_bits_pte_d ),
       .io_requestor_1_resp_bits_pte_r( ptw_io_requestor_1_resp_bits_pte_r ),
       .io_requestor_1_resp_bits_pte_typ( ptw_io_requestor_1_resp_bits_pte_typ ),
       .io_requestor_1_resp_bits_pte_v( ptw_io_requestor_1_resp_bits_pte_v ),
       .io_requestor_1_status_sd( ptw_io_requestor_1_status_sd ),
       .io_requestor_1_status_zero2( ptw_io_requestor_1_status_zero2 ),
       .io_requestor_1_status_sd_rv32( ptw_io_requestor_1_status_sd_rv32 ),
       .io_requestor_1_status_zero1( ptw_io_requestor_1_status_zero1 ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_mprv( ptw_io_requestor_1_status_mprv ),
       .io_requestor_1_status_xs( ptw_io_requestor_1_status_xs ),
       .io_requestor_1_status_fs( ptw_io_requestor_1_status_fs ),
       .io_requestor_1_status_prv3( ptw_io_requestor_1_status_prv3 ),
       .io_requestor_1_status_ie3( ptw_io_requestor_1_status_ie3 ),
       .io_requestor_1_status_prv2( ptw_io_requestor_1_status_prv2 ),
       .io_requestor_1_status_ie2( ptw_io_requestor_1_status_ie2 ),
       .io_requestor_1_status_prv1( ptw_io_requestor_1_status_prv1 ),
       .io_requestor_1_status_ie1( ptw_io_requestor_1_status_ie1 ),
       .io_requestor_1_status_prv( ptw_io_requestor_1_status_prv ),
       .io_requestor_1_status_ie( ptw_io_requestor_1_status_ie ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_ptw_req_valid ),
       .io_requestor_0_req_bits_addr( icache_io_ptw_req_bits_addr ),
       .io_requestor_0_req_bits_prv( icache_io_ptw_req_bits_prv ),
       .io_requestor_0_req_bits_store( icache_io_ptw_req_bits_store ),
       .io_requestor_0_req_bits_fetch( icache_io_ptw_req_bits_fetch ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_pte_ppn( ptw_io_requestor_0_resp_bits_pte_ppn ),
       .io_requestor_0_resp_bits_pte_reserved_for_software( ptw_io_requestor_0_resp_bits_pte_reserved_for_software ),
       .io_requestor_0_resp_bits_pte_d( ptw_io_requestor_0_resp_bits_pte_d ),
       .io_requestor_0_resp_bits_pte_r( ptw_io_requestor_0_resp_bits_pte_r ),
       .io_requestor_0_resp_bits_pte_typ( ptw_io_requestor_0_resp_bits_pte_typ ),
       .io_requestor_0_resp_bits_pte_v( ptw_io_requestor_0_resp_bits_pte_v ),
       .io_requestor_0_status_sd( ptw_io_requestor_0_status_sd ),
       .io_requestor_0_status_zero2( ptw_io_requestor_0_status_zero2 ),
       .io_requestor_0_status_sd_rv32( ptw_io_requestor_0_status_sd_rv32 ),
       .io_requestor_0_status_zero1( ptw_io_requestor_0_status_zero1 ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_mprv( ptw_io_requestor_0_status_mprv ),
       .io_requestor_0_status_xs( ptw_io_requestor_0_status_xs ),
       .io_requestor_0_status_fs( ptw_io_requestor_0_status_fs ),
       .io_requestor_0_status_prv3( ptw_io_requestor_0_status_prv3 ),
       .io_requestor_0_status_ie3( ptw_io_requestor_0_status_ie3 ),
       .io_requestor_0_status_prv2( ptw_io_requestor_0_status_prv2 ),
       .io_requestor_0_status_ie2( ptw_io_requestor_0_status_ie2 ),
       .io_requestor_0_status_prv1( ptw_io_requestor_0_status_prv1 ),
       .io_requestor_0_status_ie1( ptw_io_requestor_0_status_ie1 ),
       .io_requestor_0_status_prv( ptw_io_requestor_0_status_prv ),
       .io_requestor_0_status_ie( ptw_io_requestor_0_status_ie ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_mem_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_data( ptw_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data_word_bypass( dcArb_io_requestor_0_resp_bits_data_word_bypass ),
       .io_mem_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_invalidate_lr(  )
       .io_mem_ordered( dcArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_status_sd( core_io_ptw_status_sd ),
       .io_dpath_status_zero2( core_io_ptw_status_zero2 ),
       .io_dpath_status_sd_rv32( core_io_ptw_status_sd_rv32 ),
       .io_dpath_status_zero1( core_io_ptw_status_zero1 ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_mprv( core_io_ptw_status_mprv ),
       .io_dpath_status_xs( core_io_ptw_status_xs ),
       .io_dpath_status_fs( core_io_ptw_status_fs ),
       .io_dpath_status_prv3( core_io_ptw_status_prv3 ),
       .io_dpath_status_ie3( core_io_ptw_status_ie3 ),
       .io_dpath_status_prv2( core_io_ptw_status_prv2 ),
       .io_dpath_status_ie2( core_io_ptw_status_ie2 ),
       .io_dpath_status_prv1( core_io_ptw_status_prv1 ),
       .io_dpath_status_ie1( core_io_ptw_status_ie1 ),
       .io_dpath_status_prv( core_io_ptw_status_prv ),
       .io_dpath_status_ie( core_io_ptw_status_ie )
  );
  HellaCacheArbiter dcArb(.clk(clk),
       .io_requestor_1_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data_word_bypass( dcArb_io_requestor_1_resp_bits_data_word_bypass ),
       .io_requestor_1_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       .io_requestor_1_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_requestor_1_ordered( dcArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_data( ptw_io_mem_req_bits_data ),
       .io_requestor_0_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data_word_bypass( dcArb_io_requestor_0_resp_bits_data_word_bypass ),
       .io_requestor_0_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_invalidate_lr(  )
       .io_requestor_0_ordered( dcArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcArb_io_mem_req_valid ),
       .io_mem_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_mem_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data_word_bypass( dcache_io_cpu_resp_bits_data_word_bypass ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_invalidate_lr(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign dcArb.io_requestor_0_req_bits_tag = {1{$random}};
// synthesis translate_on
`endif
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [11:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[11:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[63:0] T10;
  wire[76:0] T11;
  reg [76:0] ram [1:0];
  wire[76:0] T12;
  wire[76:0] T13;
  wire[76:0] T14;
  wire[75:0] T15;
  wire[11:0] T16;
  wire T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[6'h3f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_rw, T15};
  assign T15 = {io_enq_bits_addr, io_enq_bits_data};
  assign io_deq_bits_addr = T16;
  assign T16 = T11[7'h4b:7'h40];
  assign io_deq_bits_rw = T17;
  assign T17 = T11[7'h4c:7'h4c];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire[63:0] T10;
  reg [63:0] ram [1:0];
  wire[63:0] T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire T10;
  reg [0:0] ram [1:0];
  wire T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module Top(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_csr,
    input  io_mem_backup_ctrl_en,
    input  io_mem_backup_ctrl_in_valid,
    input  io_mem_backup_ctrl_out_ready,
    output io_mem_backup_ctrl_out_valid,
    input  io_mem_0_aw_ready,
    output io_mem_0_aw_valid,
    output[31:0] io_mem_0_aw_bits_addr,
    output[7:0] io_mem_0_aw_bits_len,
    output[2:0] io_mem_0_aw_bits_size,
    output[1:0] io_mem_0_aw_bits_burst,
    output io_mem_0_aw_bits_lock,
    output[3:0] io_mem_0_aw_bits_cache,
    output[2:0] io_mem_0_aw_bits_prot,
    output[3:0] io_mem_0_aw_bits_qos,
    output[3:0] io_mem_0_aw_bits_region,
    output[4:0] io_mem_0_aw_bits_id,
    output io_mem_0_aw_bits_user,
    input  io_mem_0_w_ready,
    output io_mem_0_w_valid,
    output[63:0] io_mem_0_w_bits_data,
    output io_mem_0_w_bits_last,
    output[7:0] io_mem_0_w_bits_strb,
    output io_mem_0_w_bits_user,
    output io_mem_0_b_ready,
    input  io_mem_0_b_valid,
    input [1:0] io_mem_0_b_bits_resp,
    input [4:0] io_mem_0_b_bits_id,
    input  io_mem_0_b_bits_user,
    input  io_mem_0_ar_ready,
    output io_mem_0_ar_valid,
    output[31:0] io_mem_0_ar_bits_addr,
    output[7:0] io_mem_0_ar_bits_len,
    output[2:0] io_mem_0_ar_bits_size,
    output[1:0] io_mem_0_ar_bits_burst,
    output io_mem_0_ar_bits_lock,
    output[3:0] io_mem_0_ar_bits_cache,
    output[2:0] io_mem_0_ar_bits_prot,
    output[3:0] io_mem_0_ar_bits_qos,
    output[3:0] io_mem_0_ar_bits_region,
    output[4:0] io_mem_0_ar_bits_id,
    output io_mem_0_ar_bits_user,
    output io_mem_0_r_ready,
    input  io_mem_0_r_valid,
    input [1:0] io_mem_0_r_bits_resp,
    input [63:0] io_mem_0_r_bits_data,
    input  io_mem_0_r_bits_last,
    input [4:0] io_mem_0_r_bits_id,
    input  io_mem_0_r_bits_user
);

  reg  R0;
  reg  R1;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire Queue_io_deq_bits_rw;
  wire[11:0] Queue_io_deq_bits_addr;
  wire[63:0] Queue_io_deq_bits_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire Queue_2_io_deq_bits;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire Queue_3_io_deq_bits;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[31:0] Queue_4_io_deq_bits_addr;
  wire[7:0] Queue_4_io_deq_bits_len;
  wire[2:0] Queue_4_io_deq_bits_size;
  wire[1:0] Queue_4_io_deq_bits_burst;
  wire Queue_4_io_deq_bits_lock;
  wire[2:0] Queue_4_io_deq_bits_prot;
  wire[3:0] Queue_4_io_deq_bits_qos;
  wire[3:0] Queue_4_io_deq_bits_region;
  wire[4:0] Queue_4_io_deq_bits_id;
  wire Queue_4_io_deq_bits_user;
  wire Queue_5_io_enq_ready;
  wire Queue_5_io_deq_valid;
  wire[31:0] Queue_5_io_deq_bits_addr;
  wire[7:0] Queue_5_io_deq_bits_len;
  wire[2:0] Queue_5_io_deq_bits_size;
  wire[1:0] Queue_5_io_deq_bits_burst;
  wire Queue_5_io_deq_bits_lock;
  wire[2:0] Queue_5_io_deq_bits_prot;
  wire[3:0] Queue_5_io_deq_bits_qos;
  wire[3:0] Queue_5_io_deq_bits_region;
  wire[4:0] Queue_5_io_deq_bits_id;
  wire Queue_5_io_deq_bits_user;
  wire Queue_6_io_enq_ready;
  wire Queue_6_io_deq_valid;
  wire[63:0] Queue_6_io_deq_bits_data;
  wire Queue_6_io_deq_bits_last;
  wire[7:0] Queue_6_io_deq_bits_strb;
  wire Queue_6_io_deq_bits_user;
  wire Queue_7_io_enq_ready;
  wire Queue_7_io_deq_valid;
  wire[1:0] Queue_7_io_deq_bits_resp;
  wire[63:0] Queue_7_io_deq_bits_data;
  wire Queue_7_io_deq_bits_last;
  wire[4:0] Queue_7_io_deq_bits_id;
  wire Queue_7_io_deq_bits_user;
  wire Queue_8_io_enq_ready;
  wire Queue_8_io_deq_valid;
  wire[1:0] Queue_8_io_deq_bits_resp;
  wire[4:0] Queue_8_io_deq_bits_id;
  wire Queue_8_io_deq_bits_user;
  wire errslave_io_aw_ready;
  wire errslave_io_w_ready;
  wire errslave_io_b_valid;
  wire[1:0] errslave_io_b_bits_resp;
  wire[4:0] errslave_io_b_bits_id;
  wire errslave_io_ar_ready;
  wire errslave_io_r_valid;
  wire[1:0] errslave_io_r_bits_resp;
  wire[63:0] errslave_io_r_bits_data;
  wire errslave_io_r_bits_last;
  wire[4:0] errslave_io_r_bits_id;
  wire RocketTile_io_cached_0_acquire_valid;
  wire[25:0] RocketTile_io_cached_0_acquire_bits_addr_block;
  wire[1:0] RocketTile_io_cached_0_acquire_bits_client_xact_id;
  wire[1:0] RocketTile_io_cached_0_acquire_bits_addr_beat;
  wire RocketTile_io_cached_0_acquire_bits_is_builtin_type;
  wire[2:0] RocketTile_io_cached_0_acquire_bits_a_type;
  wire[16:0] RocketTile_io_cached_0_acquire_bits_union;
  wire[127:0] RocketTile_io_cached_0_acquire_bits_data;
  wire RocketTile_io_cached_0_grant_ready;
  wire RocketTile_io_cached_0_probe_ready;
  wire RocketTile_io_cached_0_release_valid;
  wire[1:0] RocketTile_io_cached_0_release_bits_addr_beat;
  wire[25:0] RocketTile_io_cached_0_release_bits_addr_block;
  wire[1:0] RocketTile_io_cached_0_release_bits_client_xact_id;
  wire[2:0] RocketTile_io_cached_0_release_bits_r_type;
  wire RocketTile_io_cached_0_release_bits_voluntary;
  wire[127:0] RocketTile_io_cached_0_release_bits_data;
  wire RocketTile_io_uncached_0_acquire_valid;
  wire[25:0] RocketTile_io_uncached_0_acquire_bits_addr_block;
  wire[1:0] RocketTile_io_uncached_0_acquire_bits_client_xact_id;
  wire[1:0] RocketTile_io_uncached_0_acquire_bits_addr_beat;
  wire RocketTile_io_uncached_0_acquire_bits_is_builtin_type;
  wire[2:0] RocketTile_io_uncached_0_acquire_bits_a_type;
  wire[16:0] RocketTile_io_uncached_0_acquire_bits_union;
  wire[127:0] RocketTile_io_uncached_0_acquire_bits_data;
  wire RocketTile_io_uncached_0_grant_ready;
  wire RocketTile_io_host_csr_req_ready;
  wire RocketTile_io_host_csr_resp_valid;
  wire[63:0] RocketTile_io_host_csr_resp_bits;
  wire RocketTile_io_host_ipi_req_valid;
  wire RocketTile_io_host_ipi_req_bits;
  wire RocketTile_io_host_ipi_rep_ready;
  wire RocketTile_io_host_debug_stats_csr;
  wire uncore_io_host_in_ready;
  wire uncore_io_host_out_valid;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_debug_stats_csr;
  wire uncore_io_mem_0_aw_valid;
  wire[31:0] uncore_io_mem_0_aw_bits_addr;
  wire[7:0] uncore_io_mem_0_aw_bits_len;
  wire[2:0] uncore_io_mem_0_aw_bits_size;
  wire[1:0] uncore_io_mem_0_aw_bits_burst;
  wire uncore_io_mem_0_aw_bits_lock;
  wire[3:0] uncore_io_mem_0_aw_bits_cache;
  wire[2:0] uncore_io_mem_0_aw_bits_prot;
  wire[3:0] uncore_io_mem_0_aw_bits_qos;
  wire[3:0] uncore_io_mem_0_aw_bits_region;
  wire[4:0] uncore_io_mem_0_aw_bits_id;
  wire uncore_io_mem_0_aw_bits_user;
  wire uncore_io_mem_0_w_valid;
  wire[63:0] uncore_io_mem_0_w_bits_data;
  wire uncore_io_mem_0_w_bits_last;
  wire[7:0] uncore_io_mem_0_w_bits_strb;
  wire uncore_io_mem_0_w_bits_user;
  wire uncore_io_mem_0_b_ready;
  wire uncore_io_mem_0_ar_valid;
  wire[31:0] uncore_io_mem_0_ar_bits_addr;
  wire[7:0] uncore_io_mem_0_ar_bits_len;
  wire[2:0] uncore_io_mem_0_ar_bits_size;
  wire[1:0] uncore_io_mem_0_ar_bits_burst;
  wire uncore_io_mem_0_ar_bits_lock;
  wire[3:0] uncore_io_mem_0_ar_bits_cache;
  wire[2:0] uncore_io_mem_0_ar_bits_prot;
  wire[3:0] uncore_io_mem_0_ar_bits_qos;
  wire[3:0] uncore_io_mem_0_ar_bits_region;
  wire[4:0] uncore_io_mem_0_ar_bits_id;
  wire uncore_io_mem_0_ar_bits_user;
  wire uncore_io_mem_0_r_ready;
  wire uncore_io_tiles_cached_0_acquire_ready;
  wire uncore_io_tiles_cached_0_grant_valid;
  wire[1:0] uncore_io_tiles_cached_0_grant_bits_addr_beat;
  wire[1:0] uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  wire[3:0] uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire[3:0] uncore_io_tiles_cached_0_grant_bits_g_type;
  wire[127:0] uncore_io_tiles_cached_0_grant_bits_data;
  wire uncore_io_tiles_cached_0_probe_valid;
  wire[25:0] uncore_io_tiles_cached_0_probe_bits_addr_block;
  wire[1:0] uncore_io_tiles_cached_0_probe_bits_p_type;
  wire uncore_io_tiles_cached_0_release_ready;
  wire uncore_io_tiles_uncached_0_acquire_ready;
  wire uncore_io_tiles_uncached_0_grant_valid;
  wire[1:0] uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  wire[1:0] uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire[3:0] uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire[3:0] uncore_io_tiles_uncached_0_grant_bits_g_type;
  wire[127:0] uncore_io_tiles_uncached_0_grant_bits_data;
  wire uncore_io_htif_0_reset;
  wire uncore_io_htif_0_csr_req_valid;
  wire uncore_io_htif_0_csr_req_bits_rw;
  wire[11:0] uncore_io_htif_0_csr_req_bits_addr;
  wire[63:0] uncore_io_htif_0_csr_req_bits_data;
  wire uncore_io_htif_0_csr_resp_ready;
  wire uncore_io_htif_0_ipi_req_ready;
  wire uncore_io_htif_0_ipi_rep_valid;
  wire uncore_io_htif_0_ipi_rep_bits;
  wire uncore_io_mmio_aw_valid;
  wire[31:0] uncore_io_mmio_aw_bits_addr;
  wire[7:0] uncore_io_mmio_aw_bits_len;
  wire[2:0] uncore_io_mmio_aw_bits_size;
  wire[1:0] uncore_io_mmio_aw_bits_burst;
  wire uncore_io_mmio_aw_bits_lock;
  wire[3:0] uncore_io_mmio_aw_bits_cache;
  wire[2:0] uncore_io_mmio_aw_bits_prot;
  wire[3:0] uncore_io_mmio_aw_bits_qos;
  wire[3:0] uncore_io_mmio_aw_bits_region;
  wire[4:0] uncore_io_mmio_aw_bits_id;
  wire uncore_io_mmio_aw_bits_user;
  wire uncore_io_mmio_w_valid;
  wire[63:0] uncore_io_mmio_w_bits_data;
  wire uncore_io_mmio_w_bits_last;
  wire[7:0] uncore_io_mmio_w_bits_strb;
  wire uncore_io_mmio_w_bits_user;
  wire uncore_io_mmio_b_ready;
  wire uncore_io_mmio_ar_valid;
  wire[31:0] uncore_io_mmio_ar_bits_addr;
  wire[7:0] uncore_io_mmio_ar_bits_len;
  wire[2:0] uncore_io_mmio_ar_bits_size;
  wire[1:0] uncore_io_mmio_ar_bits_burst;
  wire uncore_io_mmio_ar_bits_lock;
  wire[3:0] uncore_io_mmio_ar_bits_cache;
  wire[2:0] uncore_io_mmio_ar_bits_prot;
  wire[3:0] uncore_io_mmio_ar_bits_qos;
  wire[3:0] uncore_io_mmio_ar_bits_region;
  wire[4:0] uncore_io_mmio_ar_bits_id;
  wire uncore_io_mmio_ar_bits_user;
  wire uncore_io_mmio_r_ready;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_backup_ctrl_out_valid = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_0_r_ready = Queue_7_io_enq_ready;
  assign io_mem_0_ar_bits_user = Queue_4_io_deq_bits_user;
  assign io_mem_0_ar_bits_id = Queue_4_io_deq_bits_id;
  assign io_mem_0_ar_bits_region = Queue_4_io_deq_bits_region;
  assign io_mem_0_ar_bits_qos = Queue_4_io_deq_bits_qos;
  assign io_mem_0_ar_bits_prot = Queue_4_io_deq_bits_prot;
  assign io_mem_0_ar_bits_cache = 4'h3;
  assign io_mem_0_ar_bits_lock = Queue_4_io_deq_bits_lock;
  assign io_mem_0_ar_bits_burst = Queue_4_io_deq_bits_burst;
  assign io_mem_0_ar_bits_size = Queue_4_io_deq_bits_size;
  assign io_mem_0_ar_bits_len = Queue_4_io_deq_bits_len;
  assign io_mem_0_ar_bits_addr = Queue_4_io_deq_bits_addr;
  assign io_mem_0_ar_valid = Queue_4_io_deq_valid;
  assign io_mem_0_b_ready = Queue_8_io_enq_ready;
  assign io_mem_0_w_bits_user = Queue_6_io_deq_bits_user;
  assign io_mem_0_w_bits_strb = Queue_6_io_deq_bits_strb;
  assign io_mem_0_w_bits_last = Queue_6_io_deq_bits_last;
  assign io_mem_0_w_bits_data = Queue_6_io_deq_bits_data;
  assign io_mem_0_w_valid = Queue_6_io_deq_valid;
  assign io_mem_0_aw_bits_user = Queue_5_io_deq_bits_user;
  assign io_mem_0_aw_bits_id = Queue_5_io_deq_bits_id;
  assign io_mem_0_aw_bits_region = Queue_5_io_deq_bits_region;
  assign io_mem_0_aw_bits_qos = Queue_5_io_deq_bits_qos;
  assign io_mem_0_aw_bits_prot = Queue_5_io_deq_bits_prot;
  assign io_mem_0_aw_bits_cache = 4'h3;
  assign io_mem_0_aw_bits_lock = Queue_5_io_deq_bits_lock;
  assign io_mem_0_aw_bits_burst = Queue_5_io_deq_bits_burst;
  assign io_mem_0_aw_bits_size = Queue_5_io_deq_bits_size;
  assign io_mem_0_aw_bits_len = Queue_5_io_deq_bits_len;
  assign io_mem_0_aw_bits_addr = Queue_5_io_deq_bits_addr;
  assign io_mem_0_aw_valid = Queue_5_io_deq_valid;
  assign io_host_debug_stats_csr = uncore_io_host_debug_stats_csr;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
  Uncore uncore(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       .io_host_debug_stats_csr( uncore_io_host_debug_stats_csr ),
       .io_mem_0_aw_ready( Queue_5_io_enq_ready ),
       .io_mem_0_aw_valid( uncore_io_mem_0_aw_valid ),
       .io_mem_0_aw_bits_addr( uncore_io_mem_0_aw_bits_addr ),
       .io_mem_0_aw_bits_len( uncore_io_mem_0_aw_bits_len ),
       .io_mem_0_aw_bits_size( uncore_io_mem_0_aw_bits_size ),
       .io_mem_0_aw_bits_burst( uncore_io_mem_0_aw_bits_burst ),
       .io_mem_0_aw_bits_lock( uncore_io_mem_0_aw_bits_lock ),
       .io_mem_0_aw_bits_cache( uncore_io_mem_0_aw_bits_cache ),
       .io_mem_0_aw_bits_prot( uncore_io_mem_0_aw_bits_prot ),
       .io_mem_0_aw_bits_qos( uncore_io_mem_0_aw_bits_qos ),
       .io_mem_0_aw_bits_region( uncore_io_mem_0_aw_bits_region ),
       .io_mem_0_aw_bits_id( uncore_io_mem_0_aw_bits_id ),
       .io_mem_0_aw_bits_user( uncore_io_mem_0_aw_bits_user ),
       .io_mem_0_w_ready( Queue_6_io_enq_ready ),
       .io_mem_0_w_valid( uncore_io_mem_0_w_valid ),
       .io_mem_0_w_bits_data( uncore_io_mem_0_w_bits_data ),
       .io_mem_0_w_bits_last( uncore_io_mem_0_w_bits_last ),
       .io_mem_0_w_bits_strb( uncore_io_mem_0_w_bits_strb ),
       .io_mem_0_w_bits_user( uncore_io_mem_0_w_bits_user ),
       .io_mem_0_b_ready( uncore_io_mem_0_b_ready ),
       .io_mem_0_b_valid( Queue_8_io_deq_valid ),
       .io_mem_0_b_bits_resp( Queue_8_io_deq_bits_resp ),
       .io_mem_0_b_bits_id( Queue_8_io_deq_bits_id ),
       .io_mem_0_b_bits_user( Queue_8_io_deq_bits_user ),
       .io_mem_0_ar_ready( Queue_4_io_enq_ready ),
       .io_mem_0_ar_valid( uncore_io_mem_0_ar_valid ),
       .io_mem_0_ar_bits_addr( uncore_io_mem_0_ar_bits_addr ),
       .io_mem_0_ar_bits_len( uncore_io_mem_0_ar_bits_len ),
       .io_mem_0_ar_bits_size( uncore_io_mem_0_ar_bits_size ),
       .io_mem_0_ar_bits_burst( uncore_io_mem_0_ar_bits_burst ),
       .io_mem_0_ar_bits_lock( uncore_io_mem_0_ar_bits_lock ),
       .io_mem_0_ar_bits_cache( uncore_io_mem_0_ar_bits_cache ),
       .io_mem_0_ar_bits_prot( uncore_io_mem_0_ar_bits_prot ),
       .io_mem_0_ar_bits_qos( uncore_io_mem_0_ar_bits_qos ),
       .io_mem_0_ar_bits_region( uncore_io_mem_0_ar_bits_region ),
       .io_mem_0_ar_bits_id( uncore_io_mem_0_ar_bits_id ),
       .io_mem_0_ar_bits_user( uncore_io_mem_0_ar_bits_user ),
       .io_mem_0_r_ready( uncore_io_mem_0_r_ready ),
       .io_mem_0_r_valid( Queue_7_io_deq_valid ),
       .io_mem_0_r_bits_resp( Queue_7_io_deq_bits_resp ),
       .io_mem_0_r_bits_data( Queue_7_io_deq_bits_data ),
       .io_mem_0_r_bits_last( Queue_7_io_deq_bits_last ),
       .io_mem_0_r_bits_id( Queue_7_io_deq_bits_id ),
       .io_mem_0_r_bits_user( Queue_7_io_deq_bits_user ),
       .io_tiles_cached_0_acquire_ready( uncore_io_tiles_cached_0_acquire_ready ),
       .io_tiles_cached_0_acquire_valid( RocketTile_io_cached_0_acquire_valid ),
       .io_tiles_cached_0_acquire_bits_addr_block( RocketTile_io_cached_0_acquire_bits_addr_block ),
       .io_tiles_cached_0_acquire_bits_client_xact_id( RocketTile_io_cached_0_acquire_bits_client_xact_id ),
       .io_tiles_cached_0_acquire_bits_addr_beat( RocketTile_io_cached_0_acquire_bits_addr_beat ),
       .io_tiles_cached_0_acquire_bits_is_builtin_type( RocketTile_io_cached_0_acquire_bits_is_builtin_type ),
       .io_tiles_cached_0_acquire_bits_a_type( RocketTile_io_cached_0_acquire_bits_a_type ),
       .io_tiles_cached_0_acquire_bits_union( RocketTile_io_cached_0_acquire_bits_union ),
       .io_tiles_cached_0_acquire_bits_data( RocketTile_io_cached_0_acquire_bits_data ),
       .io_tiles_cached_0_grant_ready( RocketTile_io_cached_0_grant_ready ),
       .io_tiles_cached_0_grant_valid( uncore_io_tiles_cached_0_grant_valid ),
       .io_tiles_cached_0_grant_bits_addr_beat( uncore_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_tiles_cached_0_grant_bits_client_xact_id( uncore_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_tiles_cached_0_grant_bits_manager_xact_id( uncore_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_tiles_cached_0_grant_bits_is_builtin_type( uncore_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_tiles_cached_0_grant_bits_g_type( uncore_io_tiles_cached_0_grant_bits_g_type ),
       .io_tiles_cached_0_grant_bits_data( uncore_io_tiles_cached_0_grant_bits_data ),
       .io_tiles_cached_0_probe_ready( RocketTile_io_cached_0_probe_ready ),
       .io_tiles_cached_0_probe_valid( uncore_io_tiles_cached_0_probe_valid ),
       .io_tiles_cached_0_probe_bits_addr_block( uncore_io_tiles_cached_0_probe_bits_addr_block ),
       .io_tiles_cached_0_probe_bits_p_type( uncore_io_tiles_cached_0_probe_bits_p_type ),
       .io_tiles_cached_0_release_ready( uncore_io_tiles_cached_0_release_ready ),
       .io_tiles_cached_0_release_valid( RocketTile_io_cached_0_release_valid ),
       .io_tiles_cached_0_release_bits_addr_beat( RocketTile_io_cached_0_release_bits_addr_beat ),
       .io_tiles_cached_0_release_bits_addr_block( RocketTile_io_cached_0_release_bits_addr_block ),
       .io_tiles_cached_0_release_bits_client_xact_id( RocketTile_io_cached_0_release_bits_client_xact_id ),
       .io_tiles_cached_0_release_bits_r_type( RocketTile_io_cached_0_release_bits_r_type ),
       .io_tiles_cached_0_release_bits_voluntary( RocketTile_io_cached_0_release_bits_voluntary ),
       .io_tiles_cached_0_release_bits_data( RocketTile_io_cached_0_release_bits_data ),
       .io_tiles_uncached_0_acquire_ready( uncore_io_tiles_uncached_0_acquire_ready ),
       .io_tiles_uncached_0_acquire_valid( RocketTile_io_uncached_0_acquire_valid ),
       .io_tiles_uncached_0_acquire_bits_addr_block( RocketTile_io_uncached_0_acquire_bits_addr_block ),
       .io_tiles_uncached_0_acquire_bits_client_xact_id( RocketTile_io_uncached_0_acquire_bits_client_xact_id ),
       .io_tiles_uncached_0_acquire_bits_addr_beat( RocketTile_io_uncached_0_acquire_bits_addr_beat ),
       .io_tiles_uncached_0_acquire_bits_is_builtin_type( RocketTile_io_uncached_0_acquire_bits_is_builtin_type ),
       .io_tiles_uncached_0_acquire_bits_a_type( RocketTile_io_uncached_0_acquire_bits_a_type ),
       .io_tiles_uncached_0_acquire_bits_union( RocketTile_io_uncached_0_acquire_bits_union ),
       .io_tiles_uncached_0_acquire_bits_data( RocketTile_io_uncached_0_acquire_bits_data ),
       .io_tiles_uncached_0_grant_ready( RocketTile_io_uncached_0_grant_ready ),
       .io_tiles_uncached_0_grant_valid( uncore_io_tiles_uncached_0_grant_valid ),
       .io_tiles_uncached_0_grant_bits_addr_beat( uncore_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_tiles_uncached_0_grant_bits_client_xact_id( uncore_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_tiles_uncached_0_grant_bits_manager_xact_id( uncore_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_tiles_uncached_0_grant_bits_is_builtin_type( uncore_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_tiles_uncached_0_grant_bits_g_type( uncore_io_tiles_uncached_0_grant_bits_g_type ),
       .io_tiles_uncached_0_grant_bits_data( uncore_io_tiles_uncached_0_grant_bits_data ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_csr_req_ready( Queue_io_enq_ready ),
       .io_htif_0_csr_req_valid( uncore_io_htif_0_csr_req_valid ),
       .io_htif_0_csr_req_bits_rw( uncore_io_htif_0_csr_req_bits_rw ),
       .io_htif_0_csr_req_bits_addr( uncore_io_htif_0_csr_req_bits_addr ),
       .io_htif_0_csr_req_bits_data( uncore_io_htif_0_csr_req_bits_data ),
       .io_htif_0_csr_resp_ready( uncore_io_htif_0_csr_resp_ready ),
       .io_htif_0_csr_resp_valid( Queue_1_io_deq_valid ),
       .io_htif_0_csr_resp_bits( Queue_1_io_deq_bits ),
       .io_htif_0_ipi_req_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_htif_0_ipi_req_valid( Queue_2_io_deq_valid ),
       .io_htif_0_ipi_req_bits( Queue_2_io_deq_bits ),
       .io_htif_0_ipi_rep_ready( Queue_3_io_enq_ready ),
       .io_htif_0_ipi_rep_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_htif_0_ipi_rep_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_htif_0_debug_stats_csr( RocketTile_io_host_debug_stats_csr ),
       //.io_mem_backup_ctrl_en(  )
       //.io_mem_backup_ctrl_in_valid(  )
       //.io_mem_backup_ctrl_out_ready(  )
       //.io_mem_backup_ctrl_out_valid(  )
       .io_mmio_aw_ready( errslave_io_aw_ready ),
       .io_mmio_aw_valid( uncore_io_mmio_aw_valid ),
       .io_mmio_aw_bits_addr( uncore_io_mmio_aw_bits_addr ),
       .io_mmio_aw_bits_len( uncore_io_mmio_aw_bits_len ),
       .io_mmio_aw_bits_size( uncore_io_mmio_aw_bits_size ),
       .io_mmio_aw_bits_burst( uncore_io_mmio_aw_bits_burst ),
       .io_mmio_aw_bits_lock( uncore_io_mmio_aw_bits_lock ),
       .io_mmio_aw_bits_cache( uncore_io_mmio_aw_bits_cache ),
       .io_mmio_aw_bits_prot( uncore_io_mmio_aw_bits_prot ),
       .io_mmio_aw_bits_qos( uncore_io_mmio_aw_bits_qos ),
       .io_mmio_aw_bits_region( uncore_io_mmio_aw_bits_region ),
       .io_mmio_aw_bits_id( uncore_io_mmio_aw_bits_id ),
       .io_mmio_aw_bits_user( uncore_io_mmio_aw_bits_user ),
       .io_mmio_w_ready( errslave_io_w_ready ),
       .io_mmio_w_valid( uncore_io_mmio_w_valid ),
       .io_mmio_w_bits_data( uncore_io_mmio_w_bits_data ),
       .io_mmio_w_bits_last( uncore_io_mmio_w_bits_last ),
       .io_mmio_w_bits_strb( uncore_io_mmio_w_bits_strb ),
       .io_mmio_w_bits_user( uncore_io_mmio_w_bits_user ),
       .io_mmio_b_ready( uncore_io_mmio_b_ready ),
       .io_mmio_b_valid( errslave_io_b_valid ),
       .io_mmio_b_bits_resp( errslave_io_b_bits_resp ),
       .io_mmio_b_bits_id( errslave_io_b_bits_id ),
       //.io_mmio_b_bits_user(  )
       .io_mmio_ar_ready( errslave_io_ar_ready ),
       .io_mmio_ar_valid( uncore_io_mmio_ar_valid ),
       .io_mmio_ar_bits_addr( uncore_io_mmio_ar_bits_addr ),
       .io_mmio_ar_bits_len( uncore_io_mmio_ar_bits_len ),
       .io_mmio_ar_bits_size( uncore_io_mmio_ar_bits_size ),
       .io_mmio_ar_bits_burst( uncore_io_mmio_ar_bits_burst ),
       .io_mmio_ar_bits_lock( uncore_io_mmio_ar_bits_lock ),
       .io_mmio_ar_bits_cache( uncore_io_mmio_ar_bits_cache ),
       .io_mmio_ar_bits_prot( uncore_io_mmio_ar_bits_prot ),
       .io_mmio_ar_bits_qos( uncore_io_mmio_ar_bits_qos ),
       .io_mmio_ar_bits_region( uncore_io_mmio_ar_bits_region ),
       .io_mmio_ar_bits_id( uncore_io_mmio_ar_bits_id ),
       .io_mmio_ar_bits_user( uncore_io_mmio_ar_bits_user ),
       .io_mmio_r_ready( uncore_io_mmio_r_ready ),
       .io_mmio_r_valid( errslave_io_r_valid ),
       .io_mmio_r_bits_resp( errslave_io_r_bits_resp ),
       .io_mmio_r_bits_data( errslave_io_r_bits_data ),
       .io_mmio_r_bits_last( errslave_io_r_bits_last ),
       .io_mmio_r_bits_id( errslave_io_r_bits_id )
       //.io_mmio_r_bits_user(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign uncore.io_htif_0_ipi_rep_bits = {1{$random}};
    assign uncore.io_mmio_b_bits_user = {1{$random}};
    assign uncore.io_mmio_r_bits_user = {1{$random}};
// synthesis translate_on
`endif
  RocketTile RocketTile(.clk(clk), .reset(uncore_io_htif_0_reset),
       .io_cached_0_acquire_ready( uncore_io_tiles_cached_0_acquire_ready ),
       .io_cached_0_acquire_valid( RocketTile_io_cached_0_acquire_valid ),
       .io_cached_0_acquire_bits_addr_block( RocketTile_io_cached_0_acquire_bits_addr_block ),
       .io_cached_0_acquire_bits_client_xact_id( RocketTile_io_cached_0_acquire_bits_client_xact_id ),
       .io_cached_0_acquire_bits_addr_beat( RocketTile_io_cached_0_acquire_bits_addr_beat ),
       .io_cached_0_acquire_bits_is_builtin_type( RocketTile_io_cached_0_acquire_bits_is_builtin_type ),
       .io_cached_0_acquire_bits_a_type( RocketTile_io_cached_0_acquire_bits_a_type ),
       .io_cached_0_acquire_bits_union( RocketTile_io_cached_0_acquire_bits_union ),
       .io_cached_0_acquire_bits_data( RocketTile_io_cached_0_acquire_bits_data ),
       .io_cached_0_grant_ready( RocketTile_io_cached_0_grant_ready ),
       .io_cached_0_grant_valid( uncore_io_tiles_cached_0_grant_valid ),
       .io_cached_0_grant_bits_addr_beat( uncore_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_cached_0_grant_bits_client_xact_id( uncore_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_cached_0_grant_bits_manager_xact_id( uncore_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_cached_0_grant_bits_is_builtin_type( uncore_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_cached_0_grant_bits_g_type( uncore_io_tiles_cached_0_grant_bits_g_type ),
       .io_cached_0_grant_bits_data( uncore_io_tiles_cached_0_grant_bits_data ),
       .io_cached_0_probe_ready( RocketTile_io_cached_0_probe_ready ),
       .io_cached_0_probe_valid( uncore_io_tiles_cached_0_probe_valid ),
       .io_cached_0_probe_bits_addr_block( uncore_io_tiles_cached_0_probe_bits_addr_block ),
       .io_cached_0_probe_bits_p_type( uncore_io_tiles_cached_0_probe_bits_p_type ),
       .io_cached_0_release_ready( uncore_io_tiles_cached_0_release_ready ),
       .io_cached_0_release_valid( RocketTile_io_cached_0_release_valid ),
       .io_cached_0_release_bits_addr_beat( RocketTile_io_cached_0_release_bits_addr_beat ),
       .io_cached_0_release_bits_addr_block( RocketTile_io_cached_0_release_bits_addr_block ),
       .io_cached_0_release_bits_client_xact_id( RocketTile_io_cached_0_release_bits_client_xact_id ),
       .io_cached_0_release_bits_r_type( RocketTile_io_cached_0_release_bits_r_type ),
       .io_cached_0_release_bits_voluntary( RocketTile_io_cached_0_release_bits_voluntary ),
       .io_cached_0_release_bits_data( RocketTile_io_cached_0_release_bits_data ),
       .io_uncached_0_acquire_ready( uncore_io_tiles_uncached_0_acquire_ready ),
       .io_uncached_0_acquire_valid( RocketTile_io_uncached_0_acquire_valid ),
       .io_uncached_0_acquire_bits_addr_block( RocketTile_io_uncached_0_acquire_bits_addr_block ),
       .io_uncached_0_acquire_bits_client_xact_id( RocketTile_io_uncached_0_acquire_bits_client_xact_id ),
       .io_uncached_0_acquire_bits_addr_beat( RocketTile_io_uncached_0_acquire_bits_addr_beat ),
       .io_uncached_0_acquire_bits_is_builtin_type( RocketTile_io_uncached_0_acquire_bits_is_builtin_type ),
       .io_uncached_0_acquire_bits_a_type( RocketTile_io_uncached_0_acquire_bits_a_type ),
       .io_uncached_0_acquire_bits_union( RocketTile_io_uncached_0_acquire_bits_union ),
       .io_uncached_0_acquire_bits_data( RocketTile_io_uncached_0_acquire_bits_data ),
       .io_uncached_0_grant_ready( RocketTile_io_uncached_0_grant_ready ),
       .io_uncached_0_grant_valid( uncore_io_tiles_uncached_0_grant_valid ),
       .io_uncached_0_grant_bits_addr_beat( uncore_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_uncached_0_grant_bits_client_xact_id( uncore_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_uncached_0_grant_bits_manager_xact_id( uncore_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_uncached_0_grant_bits_is_builtin_type( uncore_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_uncached_0_grant_bits_g_type( uncore_io_tiles_uncached_0_grant_bits_g_type ),
       .io_uncached_0_grant_bits_data( uncore_io_tiles_uncached_0_grant_bits_data ),
       .io_host_reset( R0 ),
       .io_host_id( 1'h0 ),
       .io_host_csr_req_ready( RocketTile_io_host_csr_req_ready ),
       .io_host_csr_req_valid( Queue_io_deq_valid ),
       .io_host_csr_req_bits_rw( Queue_io_deq_bits_rw ),
       .io_host_csr_req_bits_addr( Queue_io_deq_bits_addr ),
       .io_host_csr_req_bits_data( Queue_io_deq_bits_data ),
       .io_host_csr_resp_ready( Queue_1_io_enq_ready ),
       .io_host_csr_resp_valid( RocketTile_io_host_csr_resp_valid ),
       .io_host_csr_resp_bits( RocketTile_io_host_csr_resp_bits ),
       .io_host_ipi_req_ready( Queue_2_io_enq_ready ),
       .io_host_ipi_req_valid( RocketTile_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( RocketTile_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( RocketTile_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( Queue_3_io_deq_valid ),
       .io_host_ipi_rep_bits( Queue_3_io_deq_bits ),
       .io_host_debug_stats_csr( RocketTile_io_host_debug_stats_csr )
  );
  Queue_0 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_csr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_csr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_csr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_csr_req_bits_data ),
       .io_deq_ready( RocketTile_io_host_csr_req_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_rw( Queue_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_io_deq_bits_data )
       //.io_count(  )
  );
  Queue_1 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_csr_resp_valid ),
       .io_enq_bits( RocketTile_io_host_csr_resp_bits ),
       .io_deq_ready( uncore_io_htif_0_csr_resp_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
       //.io_count(  )
  );
  Queue_2 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_ipi_req_valid ),
       .io_enq_bits( RocketTile_io_host_ipi_req_bits ),
       .io_deq_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits( Queue_2_io_deq_bits )
       //.io_count(  )
  );
  Queue_2 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_enq_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_deq_ready( RocketTile_io_host_ipi_rep_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits( Queue_3_io_deq_bits )
       //.io_count(  )
  );
  Queue_3 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( uncore_io_mem_0_ar_valid ),
       .io_enq_bits_addr( uncore_io_mem_0_ar_bits_addr ),
       .io_enq_bits_len( uncore_io_mem_0_ar_bits_len ),
       .io_enq_bits_size( uncore_io_mem_0_ar_bits_size ),
       .io_enq_bits_burst( uncore_io_mem_0_ar_bits_burst ),
       .io_enq_bits_lock( uncore_io_mem_0_ar_bits_lock ),
       .io_enq_bits_cache( uncore_io_mem_0_ar_bits_cache ),
       .io_enq_bits_prot( uncore_io_mem_0_ar_bits_prot ),
       .io_enq_bits_qos( uncore_io_mem_0_ar_bits_qos ),
       .io_enq_bits_region( uncore_io_mem_0_ar_bits_region ),
       .io_enq_bits_id( uncore_io_mem_0_ar_bits_id ),
       .io_enq_bits_user( uncore_io_mem_0_ar_bits_user ),
       .io_deq_ready( io_mem_0_ar_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_addr( Queue_4_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_4_io_deq_bits_len ),
       .io_deq_bits_size( Queue_4_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_4_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_4_io_deq_bits_lock ),
       //.io_deq_bits_cache(  )
       .io_deq_bits_prot( Queue_4_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_4_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_4_io_deq_bits_region ),
       .io_deq_bits_id( Queue_4_io_deq_bits_id ),
       .io_deq_bits_user( Queue_4_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_3 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( uncore_io_mem_0_aw_valid ),
       .io_enq_bits_addr( uncore_io_mem_0_aw_bits_addr ),
       .io_enq_bits_len( uncore_io_mem_0_aw_bits_len ),
       .io_enq_bits_size( uncore_io_mem_0_aw_bits_size ),
       .io_enq_bits_burst( uncore_io_mem_0_aw_bits_burst ),
       .io_enq_bits_lock( uncore_io_mem_0_aw_bits_lock ),
       .io_enq_bits_cache( uncore_io_mem_0_aw_bits_cache ),
       .io_enq_bits_prot( uncore_io_mem_0_aw_bits_prot ),
       .io_enq_bits_qos( uncore_io_mem_0_aw_bits_qos ),
       .io_enq_bits_region( uncore_io_mem_0_aw_bits_region ),
       .io_enq_bits_id( uncore_io_mem_0_aw_bits_id ),
       .io_enq_bits_user( uncore_io_mem_0_aw_bits_user ),
       .io_deq_ready( io_mem_0_aw_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_addr( Queue_5_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_5_io_deq_bits_len ),
       .io_deq_bits_size( Queue_5_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_5_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_5_io_deq_bits_lock ),
       //.io_deq_bits_cache(  )
       .io_deq_bits_prot( Queue_5_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_5_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_5_io_deq_bits_region ),
       .io_deq_bits_id( Queue_5_io_deq_bits_id ),
       .io_deq_bits_user( Queue_5_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_4 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( uncore_io_mem_0_w_valid ),
       .io_enq_bits_data( uncore_io_mem_0_w_bits_data ),
       .io_enq_bits_last( uncore_io_mem_0_w_bits_last ),
       .io_enq_bits_strb( uncore_io_mem_0_w_bits_strb ),
       .io_enq_bits_user( uncore_io_mem_0_w_bits_user ),
       .io_deq_ready( io_mem_0_w_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_data( Queue_6_io_deq_bits_data ),
       .io_deq_bits_last( Queue_6_io_deq_bits_last ),
       .io_deq_bits_strb( Queue_6_io_deq_bits_strb ),
       .io_deq_bits_user( Queue_6_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_5 Queue_7(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_7_io_enq_ready ),
       .io_enq_valid( io_mem_0_r_valid ),
       .io_enq_bits_resp( io_mem_0_r_bits_resp ),
       .io_enq_bits_data( io_mem_0_r_bits_data ),
       .io_enq_bits_last( io_mem_0_r_bits_last ),
       .io_enq_bits_id( io_mem_0_r_bits_id ),
       .io_enq_bits_user( io_mem_0_r_bits_user ),
       .io_deq_ready( uncore_io_mem_0_r_ready ),
       .io_deq_valid( Queue_7_io_deq_valid ),
       .io_deq_bits_resp( Queue_7_io_deq_bits_resp ),
       .io_deq_bits_data( Queue_7_io_deq_bits_data ),
       .io_deq_bits_last( Queue_7_io_deq_bits_last ),
       .io_deq_bits_id( Queue_7_io_deq_bits_id ),
       .io_deq_bits_user( Queue_7_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_6 Queue_8(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_8_io_enq_ready ),
       .io_enq_valid( io_mem_0_b_valid ),
       .io_enq_bits_resp( io_mem_0_b_bits_resp ),
       .io_enq_bits_id( io_mem_0_b_bits_id ),
       .io_enq_bits_user( io_mem_0_b_bits_user ),
       .io_deq_ready( uncore_io_mem_0_b_ready ),
       .io_deq_valid( Queue_8_io_deq_valid ),
       .io_deq_bits_resp( Queue_8_io_deq_bits_resp ),
       .io_deq_bits_id( Queue_8_io_deq_bits_id ),
       .io_deq_bits_user( Queue_8_io_deq_bits_user )
       //.io_count(  )
  );
  NastiErrorSlave errslave(.clk(clk), .reset(reset),
       .io_aw_ready( errslave_io_aw_ready ),
       .io_aw_valid( uncore_io_mmio_aw_valid ),
       .io_aw_bits_addr( uncore_io_mmio_aw_bits_addr ),
       .io_aw_bits_len( uncore_io_mmio_aw_bits_len ),
       .io_aw_bits_size( uncore_io_mmio_aw_bits_size ),
       .io_aw_bits_burst( uncore_io_mmio_aw_bits_burst ),
       .io_aw_bits_lock( uncore_io_mmio_aw_bits_lock ),
       .io_aw_bits_cache( uncore_io_mmio_aw_bits_cache ),
       .io_aw_bits_prot( uncore_io_mmio_aw_bits_prot ),
       .io_aw_bits_qos( uncore_io_mmio_aw_bits_qos ),
       .io_aw_bits_region( uncore_io_mmio_aw_bits_region ),
       .io_aw_bits_id( uncore_io_mmio_aw_bits_id ),
       .io_aw_bits_user( uncore_io_mmio_aw_bits_user ),
       .io_w_ready( errslave_io_w_ready ),
       .io_w_valid( uncore_io_mmio_w_valid ),
       .io_w_bits_data( uncore_io_mmio_w_bits_data ),
       .io_w_bits_last( uncore_io_mmio_w_bits_last ),
       .io_w_bits_strb( uncore_io_mmio_w_bits_strb ),
       .io_w_bits_user( uncore_io_mmio_w_bits_user ),
       .io_b_ready( uncore_io_mmio_b_ready ),
       .io_b_valid( errslave_io_b_valid ),
       .io_b_bits_resp( errslave_io_b_bits_resp ),
       .io_b_bits_id( errslave_io_b_bits_id ),
       //.io_b_bits_user(  )
       .io_ar_ready( errslave_io_ar_ready ),
       .io_ar_valid( uncore_io_mmio_ar_valid ),
       .io_ar_bits_addr( uncore_io_mmio_ar_bits_addr ),
       .io_ar_bits_len( uncore_io_mmio_ar_bits_len ),
       .io_ar_bits_size( uncore_io_mmio_ar_bits_size ),
       .io_ar_bits_burst( uncore_io_mmio_ar_bits_burst ),
       .io_ar_bits_lock( uncore_io_mmio_ar_bits_lock ),
       .io_ar_bits_cache( uncore_io_mmio_ar_bits_cache ),
       .io_ar_bits_prot( uncore_io_mmio_ar_bits_prot ),
       .io_ar_bits_qos( uncore_io_mmio_ar_bits_qos ),
       .io_ar_bits_region( uncore_io_mmio_ar_bits_region ),
       .io_ar_bits_id( uncore_io_mmio_ar_bits_id ),
       .io_ar_bits_user( uncore_io_mmio_ar_bits_user ),
       .io_r_ready( uncore_io_mmio_r_ready ),
       .io_r_valid( errslave_io_r_valid ),
       .io_r_bits_resp( errslave_io_r_bits_resp ),
       .io_r_bits_data( errslave_io_r_bits_data ),
       .io_r_bits_last( errslave_io_r_bits_last ),
       .io_r_bits_id( errslave_io_r_bits_id )
       //.io_r_bits_user(  )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= uncore_io_htif_0_reset;
  end
endmodule

module DataArray_T9(
  input CLK,
  input RST,
  input init,
  input [7:0] W0A,
  input W0E,
  input [127:0] W0I,
  input [127:0] W0M,
  input [7:0] R1A,
  input R1E,
  output [127:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+64) begin
    for (j=1; j<64; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][63:0] <= W0I[63:0];
  if (W0E && W0M[64]) ram[W0A][127:64] <= W0I[127:64];
end
assign R1O = ram[reg_R1A];

endmodule


module MetadataArray_tag_arr(
  input CLK,
  input RST,
  input init,
  input [5:0] W0A,
  input W0E,
  input [87:0] W0I,
  input [87:0] W0M,
  input [5:0] R1A,
  input R1E,
  output [87:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<4; i=i+22) begin
    for (j=1; j<22; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [87:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
    end
  `endif
  reg [5:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][21:0] <= W0I[21:0];
  if (W0E && W0M[22]) ram[W0A][43:22] <= W0I[43:22];
  if (W0E && W0M[44]) ram[W0A][65:44] <= W0I[65:44];
  if (W0E && W0M[66]) ram[W0A][87:66] <= W0I[87:66];
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_T241(
  input CLK,
  input RST,
  input init,
  input [7:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0I,
  output [127:0] RW0O
);

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W) ram[RW0A] <= RW0I;
end
assign RW0O = ram[reg_RW0A];

endmodule


module ICache_tag_array(
  input CLK,
  input RST,
  input init,
  input [5:0] RW0A,
  input RW0E,
  input RW0W,
  input [79:0] RW0M,
  input [79:0] RW0I,
  output [79:0] RW0O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<4; i=i+20) begin
    for (j=1; j<20; j=j+1) begin
      if (RW0M[i] != RW0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [79:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
    end
  `endif
  reg [5:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W && RW0M[0]) ram[RW0A][19:0] <= RW0I[19:0];
  if (RW0E && RW0W && RW0M[20]) ram[RW0A][39:20] <= RW0I[39:20];
  if (RW0E && RW0W && RW0M[40]) ram[RW0A][59:40] <= RW0I[59:40];
  if (RW0E && RW0W && RW0M[60]) ram[RW0A][79:60] <= RW0I[79:60];
end
assign RW0O = ram[reg_RW0A];

endmodule


