--! @defgroup main_group RISC-V System-on-Chip VHDL IP library
--! @copydoc mainpage


--! @defgroup generic_group 1. VHDL Generic Parameters
--! @ingroup main_group
--! @details VHDL generic parameters.

--! @defgroup axi4_config_generic_group AXI4 System Bus Generic Parameters
--! @ingroup generic_group
--! @details Definition of System Bus configuraiton parameters and templates
--!          methods that should be used by any master/slave device to be 
--!          compatible with Bus Controller device.


--! @defgroup verification_group 2. RTL Verificaton
--! @ingroup main_group
--! @copydoc verification_page


--! @defgroup riscv_core_group 3. RISC-V Processor
--! @ingroup main_group
--! @copydoc riscv_core_page


--! @defgroup peripheries_group 4. Peripheries
--! @ingroup main_group
--! @copydoc peripheries_page


--! @defgroup debugger_group 5. RISC-V debugger
--! @ingroup main_group
--! @copydoc debugger_page

--! @defgroup eth_setup_group Ethernet setup
--! @ingroup debugger_group
--! @copydoc eth_link

--! @defgroup debugger_api_group SW Debugger API
--! @ingroup debugger_group
--! @copydoc sw_debugger_api_link
